
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type ALU_MSG is (R_sll, R_srl, R_sra, R_add, R_addu, R_sub, R_subu, R_and, 
   R_or, R_xor, R_seq, R_sne, R_slt, R_sgt, R_sle, R_sge, R_movi2s, R_movs2i, 
   R_movf, R_movd, R_movfp2i, R_movi2fp, R_movi2t, R_movt2i, R_sltu, R_sgtu, 
   R_sleu, R_sgeu, R_mult, R_multu, J_j, J_jal, I_beqz, I_bnez, I_bfpt, I_bfpf,
   I_addi, I_addui, I_subi, I_subui, I_andi, I_ori, I_xori, I_lhi, J_rfe, 
   J_trap, I_jr, I_jalr, I_slli, I_nop, I_srli, I_srai, I_seqi, I_snei, I_slti,
   I_sgti, I_slei, I_sgei, I_lb, I_lh, I_lw, I_lbu, I_lhu, I_lf, I_ld, I_sb, 
   I_sh, I_sw, I_sf, I_sd, I_itlb, I_sltui, I_sgtui, I_sleui, I_sgeui, nop);
attribute ENUM_ENCODING of ALU_MSG : type is 
   "0000000 0000001 0000010 0000011 0000100 0000101 0000110 0000111 0001000 0001001 0001010 0001011 0001100 0001101 0001110 0001111 0010000 0010001 0010010 0010011 0010100 0010101 0010110 0010111 0011000 0011001 0011010 0011011 0011100 0011101 0011110 0011111 0100000 0100001 0100010 0100011 0100100 0100101 0100110 0100111 0101000 0101001 0101010 0101011 0101100 0101101 0101110 0101111 0110000 0110001 0110010 0110011 0110100 0110101 0110110 0110111 0111000 0111001 0111010 0111011 0111100 0111101 0111110 0111111 1000000 1000001 1000010 1000011 1000100 1000101 1000110 1000111 1001000 1001001 1001010 1001011";
type FPU_MSG is (addf, subf, multf, divf, addd, subd, multd, divd, cvtf2d, 
   cvtf2i, cvtd2f, cvtd2i, cvti2f, cvti2d, mult, div, eqf, nef, ltf, gtf, lef, 
   gef, multu, divu, eqd, ned, ltd, gtd, led, ged, nop);
attribute ENUM_ENCODING of FPU_MSG : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111 11000 11001 11010 11011 11100 11101 11110";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_ALU_MSG(arg : in std_logic_vector( 1 to 7 )) 
               return ALU_MSG;
   function ALU_MSG_to_std_logic_vector(arg : in ALU_MSG) return 
               std_logic_vector;
   function std_logic_vector_to_FPU_MSG(arg : in std_logic_vector( 1 to 5 )) 
               return FPU_MSG;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_ALU_MSG(arg : in std_logic_vector( 1 to 7 )) 
   return ALU_MSG is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000000" => return R_sll;
         when "0000001" => return R_srl;
         when "0000010" => return R_sra;
         when "0000011" => return R_add;
         when "0000100" => return R_addu;
         when "0000101" => return R_sub;
         when "0000110" => return R_subu;
         when "0000111" => return R_and;
         when "0001000" => return R_or;
         when "0001001" => return R_xor;
         when "0001010" => return R_seq;
         when "0001011" => return R_sne;
         when "0001100" => return R_slt;
         when "0001101" => return R_sgt;
         when "0001110" => return R_sle;
         when "0001111" => return R_sge;
         when "0010000" => return R_movi2s;
         when "0010001" => return R_movs2i;
         when "0010010" => return R_movf;
         when "0010011" => return R_movd;
         when "0010100" => return R_movfp2i;
         when "0010101" => return R_movi2fp;
         when "0010110" => return R_movi2t;
         when "0010111" => return R_movt2i;
         when "0011000" => return R_sltu;
         when "0011001" => return R_sgtu;
         when "0011010" => return R_sleu;
         when "0011011" => return R_sgeu;
         when "0011100" => return R_mult;
         when "0011101" => return R_multu;
         when "0011110" => return J_j;
         when "0011111" => return J_jal;
         when "0100000" => return I_beqz;
         when "0100001" => return I_bnez;
         when "0100010" => return I_bfpt;
         when "0100011" => return I_bfpf;
         when "0100100" => return I_addi;
         when "0100101" => return I_addui;
         when "0100110" => return I_subi;
         when "0100111" => return I_subui;
         when "0101000" => return I_andi;
         when "0101001" => return I_ori;
         when "0101010" => return I_xori;
         when "0101011" => return I_lhi;
         when "0101100" => return J_rfe;
         when "0101101" => return J_trap;
         when "0101110" => return I_jr;
         when "0101111" => return I_jalr;
         when "0110000" => return I_slli;
         when "0110001" => return I_nop;
         when "0110010" => return I_srli;
         when "0110011" => return I_srai;
         when "0110100" => return I_seqi;
         when "0110101" => return I_snei;
         when "0110110" => return I_slti;
         when "0110111" => return I_sgti;
         when "0111000" => return I_slei;
         when "0111001" => return I_sgei;
         when "0111010" => return I_lb;
         when "0111011" => return I_lh;
         when "0111100" => return I_lw;
         when "0111101" => return I_lbu;
         when "0111110" => return I_lhu;
         when "0111111" => return I_lf;
         when "1000000" => return I_ld;
         when "1000001" => return I_sb;
         when "1000010" => return I_sh;
         when "1000011" => return I_sw;
         when "1000100" => return I_sf;
         when "1000101" => return I_sd;
         when "1000110" => return I_itlb;
         when "1000111" => return I_sltui;
         when "1001000" => return I_sgtui;
         when "1001001" => return I_sleui;
         when "1001010" => return I_sgeui;
         when "1001011" => return nop;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return R_sll;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function ALU_MSG_to_std_logic_vector(arg : in ALU_MSG) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when R_sll => return "0000000";
         when R_srl => return "0000001";
         when R_sra => return "0000010";
         when R_add => return "0000011";
         when R_addu => return "0000100";
         when R_sub => return "0000101";
         when R_subu => return "0000110";
         when R_and => return "0000111";
         when R_or => return "0001000";
         when R_xor => return "0001001";
         when R_seq => return "0001010";
         when R_sne => return "0001011";
         when R_slt => return "0001100";
         when R_sgt => return "0001101";
         when R_sle => return "0001110";
         when R_sge => return "0001111";
         when R_movi2s => return "0010000";
         when R_movs2i => return "0010001";
         when R_movf => return "0010010";
         when R_movd => return "0010011";
         when R_movfp2i => return "0010100";
         when R_movi2fp => return "0010101";
         when R_movi2t => return "0010110";
         when R_movt2i => return "0010111";
         when R_sltu => return "0011000";
         when R_sgtu => return "0011001";
         when R_sleu => return "0011010";
         when R_sgeu => return "0011011";
         when R_mult => return "0011100";
         when R_multu => return "0011101";
         when J_j => return "0011110";
         when J_jal => return "0011111";
         when I_beqz => return "0100000";
         when I_bnez => return "0100001";
         when I_bfpt => return "0100010";
         when I_bfpf => return "0100011";
         when I_addi => return "0100100";
         when I_addui => return "0100101";
         when I_subi => return "0100110";
         when I_subui => return "0100111";
         when I_andi => return "0101000";
         when I_ori => return "0101001";
         when I_xori => return "0101010";
         when I_lhi => return "0101011";
         when J_rfe => return "0101100";
         when J_trap => return "0101101";
         when I_jr => return "0101110";
         when I_jalr => return "0101111";
         when I_slli => return "0110000";
         when I_nop => return "0110001";
         when I_srli => return "0110010";
         when I_srai => return "0110011";
         when I_seqi => return "0110100";
         when I_snei => return "0110101";
         when I_slti => return "0110110";
         when I_sgti => return "0110111";
         when I_slei => return "0111000";
         when I_sgei => return "0111001";
         when I_lb => return "0111010";
         when I_lh => return "0111011";
         when I_lw => return "0111100";
         when I_lbu => return "0111101";
         when I_lhu => return "0111110";
         when I_lf => return "0111111";
         when I_ld => return "1000000";
         when I_sb => return "1000001";
         when I_sh => return "1000010";
         when I_sw => return "1000011";
         when I_sf => return "1000100";
         when I_sd => return "1000101";
         when I_itlb => return "1000110";
         when I_sltui => return "1000111";
         when I_sgtui => return "1001000";
         when I_sleui => return "1001001";
         when I_sgeui => return "1001010";
         when nop => return "1001011";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000000";
      end case;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_FPU_MSG(arg : in std_logic_vector( 1 to 5 )) 
   return FPU_MSG is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return addf;
         when "00001" => return subf;
         when "00010" => return multf;
         when "00011" => return divf;
         when "00100" => return addd;
         when "00101" => return subd;
         when "00110" => return multd;
         when "00111" => return divd;
         when "01000" => return cvtf2d;
         when "01001" => return cvtf2i;
         when "01010" => return cvtd2f;
         when "01011" => return cvtd2i;
         when "01100" => return cvti2f;
         when "01101" => return cvti2d;
         when "01110" => return mult;
         when "01111" => return div;
         when "10000" => return eqf;
         when "10001" => return nef;
         when "10010" => return ltf;
         when "10011" => return gtf;
         when "10100" => return lef;
         when "10101" => return gef;
         when "10110" => return multu;
         when "10111" => return divu;
         when "11000" => return eqd;
         when "11001" => return ned;
         when "11010" => return ltd;
         when "11011" => return gtd;
         when "11100" => return led;
         when "11101" => return ged;
         when "11110" => return nop;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return addf;
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_addsub_3 is

   port( A, B : in std_logic_vector (32 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (32 downto 0);  CO : out std_logic);

end ALU_N32_DW01_addsub_3;

architecture SYN_cla of ALU_N32_DW01_addsub_3 is

   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => n47, A2 => n271, ZN => n1);
   U3 : AND2_X1 port map( A1 => n254, A2 => n255, ZN => n2);
   U4 : AND3_X1 port map( A1 => n59, A2 => n60, A3 => n285, ZN => n3);
   U5 : AND2_X1 port map( A1 => n228, A2 => n229, ZN => n4);
   U6 : OAI21_X1 port map( B1 => n2, B2 => n235, A => n236, ZN => n230);
   U7 : AOI21_X1 port map( B1 => n237, B2 => n238, A => n239, ZN => n235);
   U8 : OAI21_X1 port map( B1 => n1, B2 => n240, A => n241, ZN => n237);
   U9 : NAND2_X1 port map( A1 => n244, A2 => n36, ZN => n240);
   U10 : OAI21_X1 port map( B1 => n25, B2 => n135, A => n136, ZN => n133);
   U11 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n135);
   U12 : OAI21_X1 port map( B1 => n140, B2 => n141, A => n142, ZN => n137);
   U13 : NAND2_X1 port map( A1 => n144, A2 => n146, ZN => n141);
   U14 : NOR2_X1 port map( A1 => n21, A2 => n74, ZN => n73);
   U15 : AOI21_X1 port map( B1 => n230, B2 => n231, A => n232, ZN => n220);
   U16 : OAI21_X1 port map( B1 => n4, B2 => n220, A => n221, ZN => n215);
   U17 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n121);
   U18 : NAND2_X1 port map( A1 => A(6), A2 => n277, ZN => n43);
   U19 : XNOR2_X1 port map( A => n321, B => n278, ZN => n277);
   U20 : INV_X1 port map( A => B(6), ZN => n278);
   U21 : NAND2_X1 port map( A1 => n273, A2 => n274, ZN => n48);
   U22 : INV_X1 port map( A => A(7), ZN => n274);
   U23 : NAND2_X1 port map( A1 => A(7), A2 => n313, ZN => n47);
   U24 : XNOR2_X1 port map( A => n321, B => n314, ZN => n313);
   U25 : INV_X1 port map( A => B(7), ZN => n314);
   U26 : OAI21_X1 port map( B1 => n7, B2 => n207, A => n208, ZN => n205);
   U27 : OAI21_X1 port map( B1 => n18, B2 => n103, A => n104, ZN => n102);
   U28 : AOI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => n103);
   U29 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n110, ZN => n105);
   U30 : NAND2_X1 port map( A1 => n77, A2 => n80, ZN => n81);
   U31 : OR2_X1 port map( A1 => n5, A2 => A(17), ZN => n180);
   U32 : XOR2_X1 port map( A => B(17), B => n321, Z => n5);
   U33 : INV_X1 port map( A => n321, ZN => n299);
   U34 : NAND2_X1 port map( A1 => A(0), A2 => n317, ZN => n185);
   U35 : XNOR2_X1 port map( A => n321, B => n318, ZN => n317);
   U36 : INV_X1 port map( A => B(0), ZN => n318);
   U37 : NAND2_X1 port map( A1 => n319, A2 => n320, ZN => n187);
   U38 : INV_X1 port map( A => A(0), ZN => n320);
   U39 : NAND2_X1 port map( A1 => n304, A2 => n90, ZN => n300);
   U40 : NAND2_X1 port map( A1 => n90, A2 => n187, ZN => n295);
   U41 : NAND2_X1 port map( A1 => A(9), A2 => n263, ZN => n37);
   U42 : XNOR2_X1 port map( A => n321, B => n264, ZN => n263);
   U43 : INV_X1 port map( A => B(9), ZN => n264);
   U44 : NAND2_X1 port map( A1 => n265, A2 => n266, ZN => n36);
   U45 : INV_X1 port map( A => A(9), ZN => n266);
   U46 : NAND2_X1 port map( A1 => A(11), A2 => n252, ZN => n236);
   U47 : XNOR2_X1 port map( A => n321, B => n253, ZN => n252);
   U48 : INV_X1 port map( A => B(11), ZN => n253);
   U49 : NAND2_X1 port map( A1 => n259, A2 => n260, ZN => n238);
   U50 : INV_X1 port map( A => A(10), ZN => n260);
   U51 : INV_X1 port map( A => A(11), ZN => n255);
   U52 : NAND2_X1 port map( A1 => A(12), A2 => n247, ZN => n233);
   U53 : XNOR2_X1 port map( A => n321, B => n248, ZN => n247);
   U54 : INV_X1 port map( A => B(12), ZN => n248);
   U55 : NAND2_X1 port map( A1 => n245, A2 => n246, ZN => n231);
   U56 : INV_X1 port map( A => A(12), ZN => n246);
   U57 : INV_X1 port map( A => A(13), ZN => n229);
   U58 : NAND2_X1 port map( A1 => A(13), A2 => n226, ZN => n221);
   U59 : XNOR2_X1 port map( A => n321, B => n227, ZN => n226);
   U60 : INV_X1 port map( A => B(13), ZN => n227);
   U61 : AOI21_X1 port map( B1 => n215, B2 => n216, A => n217, ZN => n207);
   U62 : NAND2_X1 port map( A1 => A(16), A2 => n209, ZN => n182);
   U63 : XNOR2_X1 port map( A => n321, B => n210, ZN => n209);
   U64 : INV_X1 port map( A => B(16), ZN => n210);
   U65 : OAI21_X1 port map( B1 => n197, B2 => n198, A => n199, ZN => n193);
   U66 : AND2_X1 port map( A1 => n77, A2 => n78, ZN => n71);
   U67 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U68 : NAND2_X1 port map( A1 => A(1), A2 => n307, ZN => n87);
   U69 : XNOR2_X1 port map( A => n321, B => n308, ZN => n307);
   U70 : INV_X1 port map( A => B(1), ZN => n308);
   U71 : NAND2_X1 port map( A1 => n302, A2 => n303, ZN => n67);
   U72 : INV_X1 port map( A => A(2), ZN => n303);
   U73 : NAND2_X1 port map( A1 => A(2), A2 => n297, ZN => n64);
   U74 : XNOR2_X1 port map( A => n321, B => n298, ZN => n297);
   U75 : INV_X1 port map( A => B(2), ZN => n298);
   U76 : NAND2_X1 port map( A1 => n293, A2 => n294, ZN => n69);
   U77 : INV_X1 port map( A => A(3), ZN => n294);
   U78 : NAND2_X1 port map( A1 => A(3), A2 => n309, ZN => n68);
   U79 : XNOR2_X1 port map( A => n321, B => n310, ZN => n309);
   U80 : INV_X1 port map( A => B(3), ZN => n310);
   U81 : NAND2_X1 port map( A1 => A(4), A2 => n283, ZN => n58);
   U82 : XNOR2_X1 port map( A => n321, B => n284, ZN => n283);
   U83 : INV_X1 port map( A => B(4), ZN => n284);
   U84 : NAND2_X1 port map( A1 => n311, A2 => n312, ZN => n59);
   U85 : INV_X1 port map( A => A(4), ZN => n312);
   U86 : NAND2_X1 port map( A1 => n68, A2 => n290, ZN => n60);
   U87 : OAI21_X1 port map( B1 => n291, B2 => n292, A => n69, ZN => n290);
   U88 : OAI21_X1 port map( B1 => n295, B2 => n296, A => n64, ZN => n292);
   U89 : AOI21_X1 port map( B1 => n87, B2 => n300, A => n301, ZN => n291);
   U90 : NAND2_X1 port map( A1 => n286, A2 => n287, ZN => n54);
   U91 : INV_X1 port map( A => A(5), ZN => n287);
   U92 : NAND2_X1 port map( A1 => A(5), A2 => n281, ZN => n52);
   U93 : XNOR2_X1 port map( A => n321, B => n282, ZN => n281);
   U94 : INV_X1 port map( A => B(5), ZN => n282);
   U95 : NAND2_X1 port map( A1 => n288, A2 => n289, ZN => n46);
   U96 : INV_X1 port map( A => A(6), ZN => n289);
   U97 : OAI21_X1 port map( B1 => n3, B2 => n272, A => n48, ZN => n271);
   U98 : OAI21_X1 port map( B1 => n275, B2 => n276, A => n43, ZN => n272);
   U99 : NOR2_X1 port map( A1 => n258, A2 => n260, ZN => n239);
   U100 : XNOR2_X1 port map( A => n321, B => B(10), ZN => n258);
   U101 : AOI21_X1 port map( B1 => n193, B2 => n174, A => n175, ZN => n188);
   U102 : OAI21_X1 port map( B1 => n12, B2 => n171, A => n172, ZN => n170);
   U103 : AOI21_X1 port map( B1 => n173, B2 => n174, A => n175, ZN => n171);
   U104 : OAI21_X1 port map( B1 => n176, B2 => n177, A => n178, ZN => n173);
   U105 : NOR2_X1 port map( A1 => n157, A2 => n139, ZN => n156);
   U106 : OAI21_X1 port map( B1 => n108, B2 => n132, A => n114, ZN => n131);
   U107 : OAI21_X1 port map( B1 => n29, B2 => n96, A => n97, ZN => n95);
   U108 : AOI21_X1 port map( B1 => n154, B2 => n138, A => n139, ZN => n149);
   U109 : NOR2_X1 port map( A1 => n107, A2 => n124, ZN => n123);
   U110 : AOI21_X1 port map( B1 => n39, B2 => n36, A => n242, ZN => n241);
   U111 : NAND2_X1 port map( A1 => A(17), A2 => n201, ZN => n199);
   U112 : XNOR2_X1 port map( A => n321, B => n202, ZN => n201);
   U113 : INV_X1 port map( A => B(17), ZN => n202);
   U114 : INV_X1 port map( A => n67, ZN => n301);
   U115 : NAND2_X1 port map( A1 => n321, A2 => n67, ZN => n296);
   U116 : NAND2_X1 port map( A1 => A(8), A2 => n267, ZN => n243);
   U117 : XNOR2_X1 port map( A => n321, B => n268, ZN => n267);
   U118 : INV_X1 port map( A => B(8), ZN => n268);
   U119 : NAND2_X1 port map( A1 => n269, A2 => n270, ZN => n244);
   U120 : INV_X1 port map( A => A(8), ZN => n270);
   U121 : AOI21_X1 port map( B1 => n279, B2 => n54, A => n280, ZN => n276);
   U122 : AND2_X1 port map( A1 => n46, A2 => n54, ZN => n285);
   U123 : OAI21_X1 port map( B1 => n1, B2 => n40, A => n243, ZN => n35);
   U124 : NAND2_X1 port map( A1 => A(14), A2 => n222, ZN => n218);
   U125 : XNOR2_X1 port map( A => n321, B => n223, ZN => n222);
   U126 : INV_X1 port map( A => B(14), ZN => n223);
   U127 : OR2_X1 port map( A1 => n6, A2 => A(14), ZN => n216);
   U128 : XOR2_X1 port map( A => B(14), B => n321, Z => n6);
   U129 : NAND2_X1 port map( A1 => A(15), A2 => n213, ZN => n208);
   U130 : XNOR2_X1 port map( A => n321, B => n214, ZN => n213);
   U131 : INV_X1 port map( A => B(15), ZN => n214);
   U132 : NOR2_X1 port map( A1 => n8, A2 => A(15), ZN => n7);
   U133 : XOR2_X1 port map( A => B(15), B => n321, Z => n8);
   U134 : OR2_X1 port map( A1 => n9, A2 => A(16), ZN => n183);
   U135 : XOR2_X1 port map( A => B(16), B => n321, Z => n9);
   U136 : AOI21_X1 port map( B1 => n179, B2 => n180, A => n181, ZN => n178);
   U137 : NAND2_X1 port map( A1 => n180, A2 => n183, ZN => n177);
   U138 : OR2_X1 port map( A1 => n10, A2 => A(18), ZN => n174);
   U139 : XOR2_X1 port map( A => B(18), B => n321, Z => n10);
   U140 : NAND2_X1 port map( A1 => A(19), A2 => n191, ZN => n172);
   U141 : XNOR2_X1 port map( A => n321, B => n192, ZN => n191);
   U142 : INV_X1 port map( A => B(19), ZN => n192);
   U143 : AND2_X1 port map( A1 => n11, A2 => A(18), ZN => n175);
   U144 : XOR2_X1 port map( A => n321, B => B(18), Z => n11);
   U145 : NOR2_X1 port map( A1 => n13, A2 => A(19), ZN => n12);
   U146 : XOR2_X1 port map( A => B(19), B => n321, Z => n13);
   U147 : NAND2_X1 port map( A1 => A(20), A2 => n168, ZN => n166);
   U148 : XNOR2_X1 port map( A => n321, B => n169, ZN => n168);
   U149 : INV_X1 port map( A => B(20), ZN => n169);
   U150 : NAND2_X1 port map( A1 => A(21), A2 => n162, ZN => n160);
   U151 : XNOR2_X1 port map( A => n321, B => n163, ZN => n162);
   U152 : INV_X1 port map( A => B(21), ZN => n163);
   U153 : OR2_X1 port map( A1 => n14, A2 => A(21), ZN => n144);
   U154 : XOR2_X1 port map( A => B(21), B => n321, Z => n14);
   U155 : OR2_X1 port map( A1 => n15, A2 => A(20), ZN => n146);
   U156 : XOR2_X1 port map( A => B(20), B => n321, Z => n15);
   U157 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n142);
   U158 : NAND2_X1 port map( A1 => A(25), A2 => n129, ZN => n127);
   U159 : XNOR2_X1 port map( A => n321, B => n130, ZN => n129);
   U160 : INV_X1 port map( A => B(25), ZN => n130);
   U161 : OR2_X1 port map( A1 => n16, A2 => A(25), ZN => n112);
   U162 : XOR2_X1 port map( A => B(25), B => n321, Z => n16);
   U163 : AOI21_X1 port map( B1 => n111, B2 => n112, A => n113, ZN => n110);
   U164 : NAND2_X1 port map( A1 => n115, A2 => n112, ZN => n109);
   U165 : NAND2_X1 port map( A1 => A(27), A2 => n119, ZN => n104);
   U166 : XNOR2_X1 port map( A => n321, B => n120, ZN => n119);
   U167 : INV_X1 port map( A => B(27), ZN => n120);
   U168 : OR2_X1 port map( A1 => n17, A2 => A(26), ZN => n106);
   U169 : XOR2_X1 port map( A => B(26), B => n321, Z => n17);
   U170 : NOR2_X1 port map( A1 => n19, A2 => A(27), ZN => n18);
   U171 : XOR2_X1 port map( A => B(27), B => n321, Z => n19);
   U172 : NAND2_X1 port map( A1 => A(30), A2 => n84, ZN => n77);
   U173 : XNOR2_X1 port map( A => n321, B => n85, ZN => n84);
   U174 : INV_X1 port map( A => B(30), ZN => n85);
   U175 : OR2_X1 port map( A1 => n20, A2 => A(30), ZN => n80);
   U176 : XOR2_X1 port map( A => B(30), B => n321, Z => n20);
   U177 : OAI21_X1 port map( B1 => n82, B2 => n31, A => n83, ZN => n79);
   U178 : NAND2_X1 port map( A1 => A(31), A2 => n75, ZN => n72);
   U179 : XNOR2_X1 port map( A => n321, B => n76, ZN => n75);
   U180 : INV_X1 port map( A => B(31), ZN => n76);
   U181 : NOR2_X1 port map( A1 => n22, A2 => A(31), ZN => n21);
   U182 : XOR2_X1 port map( A => B(31), B => n321, Z => n22);
   U183 : XNOR2_X1 port map( A => n315, B => n299, ZN => SUM(0));
   U184 : NOR2_X1 port map( A1 => n316, A2 => n304, ZN => n315);
   U185 : NAND2_X1 port map( A1 => n185, A2 => n186, ZN => n89);
   U186 : NAND2_X1 port map( A1 => n321, A2 => n187, ZN => n186);
   U187 : NAND2_X1 port map( A1 => n305, A2 => n306, ZN => n90);
   U188 : INV_X1 port map( A => A(1), ZN => n306);
   U189 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n66);
   U190 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => n88);
   U191 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => n65);
   U192 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n58, ZN => n53);
   U193 : OAI21_X1 port map( B1 => n50, B2 => n51, A => n52, ZN => n45);
   U194 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => n44);
   U195 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n34);
   U196 : OAI21_X1 port map( B1 => n261, B2 => n262, A => n37, ZN => n256);
   U197 : XNOR2_X1 port map( A => n249, B => n250, ZN => SUM(11));
   U198 : NOR2_X1 port map( A1 => n2, A2 => n251, ZN => n250);
   U199 : AOI21_X1 port map( B1 => n256, B2 => n238, A => n239, ZN => n249);
   U200 : NAND2_X1 port map( A1 => n233, A2 => n231, ZN => n234);
   U201 : NOR2_X1 port map( A1 => n4, A2 => n225, ZN => n224);
   U202 : NAND2_X1 port map( A1 => n218, A2 => n216, ZN => n219);
   U203 : NOR2_X1 port map( A1 => n7, A2 => n212, ZN => n211);
   U204 : NAND2_X1 port map( A1 => n182, A2 => n183, ZN => n206);
   U205 : OAI21_X1 port map( B1 => n204, B2 => n176, A => n182, ZN => n203);
   U206 : NOR2_X1 port map( A1 => n197, A2 => n181, ZN => n200);
   U207 : NOR2_X1 port map( A1 => n196, A2 => n175, ZN => n195);
   U208 : NOR2_X1 port map( A1 => n12, A2 => n190, ZN => n189);
   U209 : NOR2_X1 port map( A1 => n165, A2 => n143, ZN => n167);
   U210 : OAI21_X1 port map( B1 => n165, B2 => n140, A => n166, ZN => n164);
   U211 : NOR2_X1 port map( A1 => n145, A2 => n158, ZN => n161);
   U212 : OR2_X1 port map( A1 => n23, A2 => A(22), ZN => n138);
   U213 : XOR2_X1 port map( A => B(22), B => n321, Z => n23);
   U214 : OAI21_X1 port map( B1 => n158, B2 => n159, A => n160, ZN => n154);
   U215 : AND2_X1 port map( A1 => n24, A2 => A(22), ZN => n139);
   U216 : XOR2_X1 port map( A => n321, B => B(22), Z => n24);
   U217 : NAND2_X1 port map( A1 => A(23), A2 => n152, ZN => n136);
   U218 : XNOR2_X1 port map( A => n321, B => n153, ZN => n152);
   U219 : INV_X1 port map( A => B(23), ZN => n153);
   U220 : NOR2_X1 port map( A1 => n26, A2 => A(23), ZN => n25);
   U221 : XOR2_X1 port map( A => B(23), B => n321, Z => n26);
   U222 : NAND2_X1 port map( A1 => A(24), A2 => n147, ZN => n114);
   U223 : XNOR2_X1 port map( A => n321, B => n148, ZN => n147);
   U224 : INV_X1 port map( A => B(24), ZN => n148);
   U225 : OR2_X1 port map( A1 => n27, A2 => A(24), ZN => n115);
   U226 : XOR2_X1 port map( A => B(24), B => n321, Z => n27);
   U227 : AND2_X1 port map( A1 => n28, A2 => A(26), ZN => n107);
   U228 : XOR2_X1 port map( A => n321, B => B(26), Z => n28);
   U229 : XNOR2_X1 port map( A => n116, B => n117, ZN => SUM(27));
   U230 : NOR2_X1 port map( A1 => n18, A2 => n118, ZN => n117);
   U231 : AOI21_X1 port map( B1 => n121, B2 => n106, A => n107, ZN => n116);
   U232 : NAND2_X1 port map( A1 => A(28), A2 => n100, ZN => n97);
   U233 : XNOR2_X1 port map( A => n321, B => n101, ZN => n100);
   U234 : INV_X1 port map( A => B(28), ZN => n101);
   U235 : NOR2_X1 port map( A1 => n30, A2 => A(28), ZN => n29);
   U236 : XOR2_X1 port map( A => B(28), B => n321, Z => n30);
   U237 : NAND2_X1 port map( A1 => A(29), A2 => n93, ZN => n83);
   U238 : XNOR2_X1 port map( A => n321, B => n94, ZN => n93);
   U239 : INV_X1 port map( A => B(29), ZN => n94);
   U240 : NOR2_X1 port map( A1 => n32, A2 => A(29), ZN => n31);
   U241 : XOR2_X1 port map( A => B(29), B => n321, Z => n32);
   U242 : OAI21_X1 port map( B1 => n21, B2 => n71, A => n72, ZN => n70);
   U243 : XNOR2_X1 port map( A => n184, B => n89, ZN => SUM(1));
   U244 : NAND2_X1 port map( A1 => n90, A2 => n87, ZN => n184);
   U245 : XNOR2_X1 port map( A => n86, B => n66, ZN => SUM(2));
   U246 : NAND2_X1 port map( A1 => n67, A2 => n64, ZN => n86);
   U247 : XNOR2_X1 port map( A => n62, B => n63, ZN => SUM(3));
   U248 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n62);
   U249 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n63);
   U250 : XNOR2_X1 port map( A => n61, B => n60, ZN => SUM(4));
   U251 : NAND2_X1 port map( A1 => n59, A2 => n58, ZN => n61);
   U252 : NAND2_X1 port map( A1 => n54, A2 => n52, ZN => n55);
   U253 : NAND2_X1 port map( A1 => n46, A2 => n43, ZN => n49);
   U254 : XNOR2_X1 port map( A => n41, B => n42, ZN => SUM(7));
   U255 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => n41);
   U256 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => n42);
   U257 : NOR2_X1 port map( A1 => n39, A2 => n40, ZN => n38);
   U258 : XNOR2_X1 port map( A => n256, B => n33, ZN => SUM(10));
   U259 : OR2_X1 port map( A1 => n257, A2 => n239, ZN => n33);
   U260 : XNOR2_X1 port map( A => n188, B => n189, ZN => SUM(19));
   U261 : NOR2_X1 port map( A1 => n25, A2 => n151, ZN => n150);
   U262 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => n134);
   U263 : NOR2_X1 port map( A1 => n125, A2 => n113, ZN => n128);
   U264 : NOR2_X1 port map( A1 => n29, A2 => n99, ZN => n98);
   U265 : NOR2_X1 port map( A1 => n92, A2 => n31, ZN => n91);
   U266 : XNOR2_X1 port map( A => n149, B => n150, ZN => SUM(23));
   U267 : XNOR2_X1 port map( A => n34, B => n35, ZN => SUM(9));
   U268 : XNOR2_X1 port map( A => n1, B => n38, ZN => SUM(8));
   U269 : XNOR2_X1 port map( A => n49, B => n45, ZN => SUM(6));
   U270 : INV_X1 port map( A => n53, ZN => n51);
   U271 : INV_X1 port map( A => n54, ZN => n50);
   U272 : XNOR2_X1 port map( A => n55, B => n53, ZN => SUM(5));
   U273 : INV_X1 port map( A => n59, ZN => n57);
   U274 : INV_X1 port map( A => n60, ZN => n56);
   U275 : XNOR2_X1 port map( A => n70, B => n299, ZN => SUM(32));
   U276 : XNOR2_X1 port map( A => n71, B => n73, ZN => SUM(31));
   U277 : INV_X1 port map( A => n72, ZN => n74);
   U278 : XNOR2_X1 port map( A => n81, B => n79, ZN => SUM(30));
   U279 : XNOR2_X1 port map( A => n82, B => n91, ZN => SUM(29));
   U280 : INV_X1 port map( A => n83, ZN => n92);
   U281 : INV_X1 port map( A => n95, ZN => n82);
   U282 : XNOR2_X1 port map( A => n96, B => n98, ZN => SUM(28));
   U283 : INV_X1 port map( A => n97, ZN => n99);
   U284 : INV_X1 port map( A => n102, ZN => n96);
   U285 : INV_X1 port map( A => n114, ZN => n111);
   U286 : INV_X1 port map( A => n104, ZN => n118);
   U287 : XNOR2_X1 port map( A => n122, B => n123, ZN => SUM(26));
   U288 : INV_X1 port map( A => n106, ZN => n124);
   U289 : INV_X1 port map( A => n121, ZN => n122);
   U290 : XNOR2_X1 port map( A => n126, B => n128, ZN => SUM(25));
   U291 : INV_X1 port map( A => n127, ZN => n113);
   U292 : INV_X1 port map( A => n112, ZN => n125);
   U293 : INV_X1 port map( A => n131, ZN => n126);
   U294 : INV_X1 port map( A => n115, ZN => n132);
   U295 : INV_X1 port map( A => n133, ZN => n108);
   U296 : XNOR2_X1 port map( A => n134, B => n133, ZN => SUM(24));
   U297 : INV_X1 port map( A => n136, ZN => n151);
   U298 : XNOR2_X1 port map( A => n155, B => n156, ZN => SUM(22));
   U299 : INV_X1 port map( A => n138, ZN => n157);
   U300 : INV_X1 port map( A => n154, ZN => n155);
   U301 : XNOR2_X1 port map( A => n159, B => n161, ZN => SUM(21));
   U302 : INV_X1 port map( A => n144, ZN => n158);
   U303 : INV_X1 port map( A => n160, ZN => n145);
   U304 : INV_X1 port map( A => n164, ZN => n159);
   U305 : XNOR2_X1 port map( A => n140, B => n167, ZN => SUM(20));
   U306 : INV_X1 port map( A => n166, ZN => n143);
   U307 : INV_X1 port map( A => n146, ZN => n165);
   U308 : INV_X1 port map( A => n170, ZN => n140);
   U309 : INV_X1 port map( A => n182, ZN => n179);
   U310 : INV_X1 port map( A => n172, ZN => n190);
   U311 : XNOR2_X1 port map( A => n194, B => n195, ZN => SUM(18));
   U312 : INV_X1 port map( A => n174, ZN => n196);
   U313 : INV_X1 port map( A => n193, ZN => n194);
   U314 : XNOR2_X1 port map( A => n198, B => n200, ZN => SUM(17));
   U315 : INV_X1 port map( A => n199, ZN => n181);
   U316 : INV_X1 port map( A => n180, ZN => n197);
   U317 : INV_X1 port map( A => n203, ZN => n198);
   U318 : INV_X1 port map( A => n205, ZN => n176);
   U319 : INV_X1 port map( A => n183, ZN => n204);
   U320 : XNOR2_X1 port map( A => n206, B => n205, ZN => SUM(16));
   U321 : XNOR2_X1 port map( A => n207, B => n211, ZN => SUM(15));
   U322 : INV_X1 port map( A => n208, ZN => n212);
   U323 : INV_X1 port map( A => n218, ZN => n217);
   U324 : XNOR2_X1 port map( A => n219, B => n215, ZN => SUM(14));
   U325 : XNOR2_X1 port map( A => n220, B => n224, ZN => SUM(13));
   U326 : INV_X1 port map( A => n221, ZN => n225);
   U327 : XNOR2_X1 port map( A => B(13), B => n321, ZN => n228);
   U328 : INV_X1 port map( A => n233, ZN => n232);
   U329 : XNOR2_X1 port map( A => n234, B => n230, ZN => SUM(12));
   U330 : INV_X1 port map( A => n37, ZN => n242);
   U331 : INV_X1 port map( A => n243, ZN => n39);
   U332 : XNOR2_X1 port map( A => B(12), B => n321, ZN => n245);
   U333 : INV_X1 port map( A => n236, ZN => n251);
   U334 : XNOR2_X1 port map( A => B(11), B => n321, ZN => n254);
   U335 : INV_X1 port map( A => n238, ZN => n257);
   U336 : XNOR2_X1 port map( A => B(10), B => n321, ZN => n259);
   U337 : INV_X1 port map( A => n36, ZN => n262);
   U338 : XNOR2_X1 port map( A => B(9), B => n321, ZN => n265);
   U339 : INV_X1 port map( A => n35, ZN => n261);
   U340 : INV_X1 port map( A => n244, ZN => n40);
   U341 : XNOR2_X1 port map( A => B(8), B => n321, ZN => n269);
   U342 : XNOR2_X1 port map( A => B(7), B => n321, ZN => n273);
   U343 : INV_X1 port map( A => n52, ZN => n280);
   U344 : INV_X1 port map( A => n58, ZN => n279);
   U345 : INV_X1 port map( A => n46, ZN => n275);
   U346 : XNOR2_X1 port map( A => B(5), B => n321, ZN => n286);
   U347 : XNOR2_X1 port map( A => B(6), B => n321, ZN => n288);
   U348 : XNOR2_X1 port map( A => B(3), B => n321, ZN => n293);
   U349 : XNOR2_X1 port map( A => B(2), B => n321, ZN => n302);
   U350 : XNOR2_X1 port map( A => B(1), B => n321, ZN => n305);
   U351 : XNOR2_X1 port map( A => B(4), B => n321, ZN => n311);
   U352 : INV_X1 port map( A => n185, ZN => n304);
   U353 : INV_X1 port map( A => n187, ZN => n316);
   U354 : XNOR2_X1 port map( A => B(0), B => n321, ZN => n319);
   U355 : BUF_X8 port map( A => ADD_SUB, Z => n321);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N5_3 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 downto 
         0);  data_out : out std_logic_vector (4 downto 0));

end gen_reg_N5_3;

architecture SYN_behav of gen_reg_N5_3 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
      n26 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n22, B2 => n16, A => n21, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n16, A2 => data_in(0), ZN => n21);
   U4 : OAI21_X1 port map( B1 => n23, B2 => n16, A => n20, ZN => n4);
   U5 : NAND2_X1 port map( A1 => data_in(1), A2 => n16, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n24, B2 => n16, A => n19, ZN => n3);
   U7 : NAND2_X1 port map( A1 => data_in(2), A2 => n16, ZN => n19);
   U8 : OAI21_X1 port map( B1 => n25, B2 => n16, A => n18, ZN => n2);
   U9 : NAND2_X1 port map( A1 => data_in(3), A2 => n16, ZN => n18);
   U10 : OAI21_X1 port map( B1 => n26, B2 => n16, A => n17, ZN => n1);
   U11 : NAND2_X1 port map( A1 => data_in(4), A2 => n16, ZN => n17);
   U12 : CLKBUF_X1 port map( A => ld, Z => n16);
   data_out_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           data_out(4), QN => n26);
   data_out_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           data_out(3), QN => n25);
   data_out_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           data_out(2), QN => n24);
   data_out_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           data_out(1), QN => n23);
   data_out_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           data_out(0), QN => n22);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N5_2 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 downto 
         0);  data_out : out std_logic_vector (4 downto 0));

end gen_reg_N5_2;

architecture SYN_behav of gen_reg_N5_2 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
      n26 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n22, B2 => n16, A => n21, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n16, A2 => data_in(0), ZN => n21);
   U4 : OAI21_X1 port map( B1 => n23, B2 => n16, A => n20, ZN => n4);
   U5 : NAND2_X1 port map( A1 => data_in(1), A2 => n16, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n24, B2 => n16, A => n19, ZN => n3);
   U7 : NAND2_X1 port map( A1 => data_in(2), A2 => n16, ZN => n19);
   U8 : OAI21_X1 port map( B1 => n25, B2 => n16, A => n18, ZN => n2);
   U9 : NAND2_X1 port map( A1 => data_in(3), A2 => n16, ZN => n18);
   U10 : OAI21_X1 port map( B1 => n26, B2 => n16, A => n17, ZN => n1);
   U11 : NAND2_X1 port map( A1 => data_in(4), A2 => n16, ZN => n17);
   U12 : CLKBUF_X1 port map( A => ld, Z => n16);
   data_out_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           data_out(4), QN => n26);
   data_out_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           data_out(3), QN => n25);
   data_out_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           data_out(2), QN => n24);
   data_out_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           data_out(1), QN => n23);
   data_out_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           data_out(0), QN => n22);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N5_1 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 downto 
         0);  data_out : out std_logic_vector (4 downto 0));

end gen_reg_N5_1;

architecture SYN_behav of gen_reg_N5_1 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
      n26 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n22, B2 => n16, A => n21, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n16, A2 => data_in(0), ZN => n21);
   U4 : OAI21_X1 port map( B1 => n23, B2 => n16, A => n20, ZN => n4);
   U5 : NAND2_X1 port map( A1 => data_in(1), A2 => n16, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n24, B2 => n16, A => n19, ZN => n3);
   U7 : NAND2_X1 port map( A1 => data_in(2), A2 => n16, ZN => n19);
   U8 : OAI21_X1 port map( B1 => n25, B2 => n16, A => n18, ZN => n2);
   U9 : NAND2_X1 port map( A1 => data_in(3), A2 => n16, ZN => n18);
   U10 : OAI21_X1 port map( B1 => n26, B2 => n16, A => n17, ZN => n1);
   U11 : NAND2_X1 port map( A1 => data_in(4), A2 => n16, ZN => n17);
   U12 : CLKBUF_X1 port map( A => ld, Z => n16);
   data_out_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           data_out(4), QN => n26);
   data_out_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           data_out(3), QN => n25);
   data_out_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           data_out(2), QN => n24);
   data_out_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           data_out(1), QN => n23);
   data_out_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           data_out(0), QN => n22);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_7 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_7;

architecture SYN_behav of gen_reg_N32_7 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n99, n108, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n174, B2 => n99, A => n147, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n108, A2 => data_in(26), ZN => n147);
   U4 : OAI21_X1 port map( B1 => n175, B2 => n108, A => n146, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(27), A2 => n108, ZN => n146);
   U6 : OAI21_X1 port map( B1 => n176, B2 => ld, A => n145, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(28), A2 => ld, ZN => n145);
   U8 : OAI21_X1 port map( B1 => n177, B2 => n108, A => n144, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(29), A2 => n108, ZN => n144);
   U10 : OAI21_X1 port map( B1 => n178, B2 => ld, A => n143, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(30), A2 => n108, ZN => n143);
   U12 : OAI21_X1 port map( B1 => n179, B2 => ld, A => n142, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(31), A2 => n108, ZN => n142);
   U14 : OAI21_X1 port map( B1 => n148, B2 => ld, A => n141, ZN => n35);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => n99, ZN => n141);
   U16 : OAI21_X1 port map( B1 => n149, B2 => ld, A => n140, ZN => n34);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n99, ZN => n140);
   U18 : OAI21_X1 port map( B1 => n150, B2 => n108, A => n139, ZN => n33);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n108, ZN => n139);
   U20 : OAI21_X1 port map( B1 => n151, B2 => n108, A => n138, ZN => n32);
   U21 : NAND2_X1 port map( A1 => data_in(3), A2 => n99, ZN => n138);
   U22 : OAI21_X1 port map( B1 => n152, B2 => ld, A => n137, ZN => n31);
   U23 : NAND2_X1 port map( A1 => data_in(4), A2 => n99, ZN => n137);
   U24 : OAI21_X1 port map( B1 => n153, B2 => ld, A => n136, ZN => n30);
   U25 : NAND2_X1 port map( A1 => data_in(5), A2 => n99, ZN => n136);
   U26 : OAI21_X1 port map( B1 => n154, B2 => n99, A => n135, ZN => n29);
   U27 : NAND2_X1 port map( A1 => data_in(6), A2 => n99, ZN => n135);
   U28 : OAI21_X1 port map( B1 => n155, B2 => ld, A => n134, ZN => n28);
   U29 : NAND2_X1 port map( A1 => data_in(7), A2 => n99, ZN => n134);
   U30 : OAI21_X1 port map( B1 => n156, B2 => n108, A => n133, ZN => n27);
   U31 : NAND2_X1 port map( A1 => data_in(8), A2 => n108, ZN => n133);
   U32 : OAI21_X1 port map( B1 => n157, B2 => ld, A => n132, ZN => n26);
   U33 : NAND2_X1 port map( A1 => data_in(9), A2 => n99, ZN => n132);
   U34 : OAI21_X1 port map( B1 => n158, B2 => ld, A => n131, ZN => n25);
   U35 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n131);
   U36 : OAI21_X1 port map( B1 => n159, B2 => ld, A => n130, ZN => n24);
   U37 : NAND2_X1 port map( A1 => data_in(11), A2 => n99, ZN => n130);
   U38 : OAI21_X1 port map( B1 => n160, B2 => n108, A => n129, ZN => n23);
   U39 : NAND2_X1 port map( A1 => data_in(12), A2 => n99, ZN => n129);
   U40 : OAI21_X1 port map( B1 => n161, B2 => n99, A => n128, ZN => n22);
   U41 : NAND2_X1 port map( A1 => data_in(13), A2 => n108, ZN => n128);
   U42 : OAI21_X1 port map( B1 => n162, B2 => n108, A => n127, ZN => n21);
   U43 : NAND2_X1 port map( A1 => data_in(14), A2 => n108, ZN => n127);
   U44 : OAI21_X1 port map( B1 => n163, B2 => ld, A => n126, ZN => n20);
   U45 : NAND2_X1 port map( A1 => data_in(15), A2 => n99, ZN => n126);
   U46 : OAI21_X1 port map( B1 => n164, B2 => ld, A => n125, ZN => n19);
   U47 : NAND2_X1 port map( A1 => data_in(16), A2 => n108, ZN => n125);
   U48 : OAI21_X1 port map( B1 => n165, B2 => n99, A => n124, ZN => n18);
   U49 : NAND2_X1 port map( A1 => data_in(17), A2 => n99, ZN => n124);
   U50 : OAI21_X1 port map( B1 => n166, B2 => n108, A => n123, ZN => n17);
   U51 : NAND2_X1 port map( A1 => data_in(18), A2 => n99, ZN => n123);
   U52 : OAI21_X1 port map( B1 => n167, B2 => ld, A => n122, ZN => n16);
   U53 : NAND2_X1 port map( A1 => data_in(19), A2 => n99, ZN => n122);
   U54 : OAI21_X1 port map( B1 => n168, B2 => n108, A => n121, ZN => n15);
   U55 : NAND2_X1 port map( A1 => data_in(20), A2 => n108, ZN => n121);
   U56 : OAI21_X1 port map( B1 => n169, B2 => n99, A => n120, ZN => n14);
   U57 : NAND2_X1 port map( A1 => data_in(21), A2 => n108, ZN => n120);
   U58 : OAI21_X1 port map( B1 => n170, B2 => n99, A => n119, ZN => n13);
   U59 : NAND2_X1 port map( A1 => data_in(22), A2 => n108, ZN => n119);
   U60 : OAI21_X1 port map( B1 => n171, B2 => ld, A => n118, ZN => n12);
   U61 : NAND2_X1 port map( A1 => data_in(23), A2 => n108, ZN => n118);
   U62 : OAI21_X1 port map( B1 => n172, B2 => n99, A => n117, ZN => n11);
   U63 : NAND2_X1 port map( A1 => data_in(24), A2 => n108, ZN => n117);
   U64 : OAI21_X1 port map( B1 => n173, B2 => n108, A => n116, ZN => n10);
   U65 : NAND2_X1 port map( A1 => data_in(25), A2 => n99, ZN => n116);
   U72 : CLKBUF_X1 port map( A => n108, Z => n99);
   U80 : CLKBUF_X1 port map( A => ld, Z => n108);
   data_out_reg_31_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n179);
   data_out_reg_30_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n178);
   data_out_reg_29_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n177);
   data_out_reg_28_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n176);
   data_out_reg_27_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n175);
   data_out_reg_26_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n174);
   data_out_reg_25_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(25), QN => n173);
   data_out_reg_24_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(24), QN => n172);
   data_out_reg_23_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(23), QN => n171);
   data_out_reg_22_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n170);
   data_out_reg_21_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n169);
   data_out_reg_20_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n168);
   data_out_reg_19_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n167);
   data_out_reg_18_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n166);
   data_out_reg_17_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n165);
   data_out_reg_16_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n164);
   data_out_reg_15_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n163);
   data_out_reg_14_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n162);
   data_out_reg_13_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n161);
   data_out_reg_12_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n160);
   data_out_reg_11_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n159);
   data_out_reg_10_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n158);
   data_out_reg_9_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n157);
   data_out_reg_8_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n156);
   data_out_reg_7_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n155);
   data_out_reg_6_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n154);
   data_out_reg_5_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n153);
   data_out_reg_4_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n152);
   data_out_reg_3_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n151);
   data_out_reg_2_inst : DFFR_X1 port map( D => n33, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n150);
   data_out_reg_1_inst : DFFR_X1 port map( D => n34, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n149);
   data_out_reg_0_inst : DFFR_X1 port map( D => n35, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n148);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_4 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_4;

architecture SYN_behav of gen_reg_N32_4 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n101, n102, n108, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n171, B2 => n101, A => n147, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n102, A2 => data_in(23), ZN => n147);
   U4 : OAI21_X1 port map( B1 => n172, B2 => n108, A => n146, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n101, ZN => n146);
   U6 : OAI21_X1 port map( B1 => n173, B2 => n101, A => n145, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => n101, ZN => n145);
   U8 : OAI21_X1 port map( B1 => n174, B2 => n102, A => n144, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => n102, ZN => n144);
   U10 : OAI21_X1 port map( B1 => n175, B2 => n102, A => n143, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => n101, ZN => n143);
   U12 : OAI21_X1 port map( B1 => n176, B2 => n108, A => n142, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => n101, ZN => n142);
   U14 : OAI21_X1 port map( B1 => n148, B2 => n101, A => n141, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => n102, ZN => n141);
   U16 : OAI21_X1 port map( B1 => n149, B2 => n101, A => n140, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n102, ZN => n140);
   U18 : OAI21_X1 port map( B1 => n150, B2 => n108, A => n139, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n102, ZN => n139);
   U20 : OAI21_X1 port map( B1 => n177, B2 => ld, A => n138, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n108, ZN => n138);
   U22 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n137, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n101, ZN => n137);
   U24 : OAI21_X1 port map( B1 => n152, B2 => n102, A => n136, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n108, ZN => n136);
   U26 : OAI21_X1 port map( B1 => n153, B2 => n102, A => n135, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n108, ZN => n135);
   U28 : OAI21_X1 port map( B1 => n154, B2 => n102, A => n134, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n108, ZN => n134);
   U30 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n133, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n108, ZN => n133);
   U32 : OAI21_X1 port map( B1 => n156, B2 => ld, A => n132, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n108, ZN => n132);
   U34 : OAI21_X1 port map( B1 => n157, B2 => ld, A => n131, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n108, ZN => n131);
   U36 : OAI21_X1 port map( B1 => n158, B2 => n102, A => n130, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n108, ZN => n130);
   U38 : OAI21_X1 port map( B1 => n159, B2 => n101, A => n129, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n102, ZN => n129);
   U40 : OAI21_X1 port map( B1 => n160, B2 => n102, A => n128, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n102, ZN => n128);
   U42 : OAI21_X1 port map( B1 => n178, B2 => n102, A => n127, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => n102, ZN => n127);
   U44 : OAI21_X1 port map( B1 => n161, B2 => n101, A => n126, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n102, ZN => n126);
   U46 : OAI21_X1 port map( B1 => n162, B2 => n108, A => n125, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => ld, ZN => n125);
   U48 : OAI21_X1 port map( B1 => n163, B2 => n108, A => n124, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => ld, ZN => n124);
   U50 : OAI21_X1 port map( B1 => n164, B2 => n102, A => n123, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => ld, ZN => n123);
   U52 : OAI21_X1 port map( B1 => n165, B2 => n102, A => n122, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n101, ZN => n122);
   U54 : OAI21_X1 port map( B1 => n166, B2 => n101, A => n121, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => ld, ZN => n121);
   U56 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n120, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n101, ZN => n120);
   U58 : OAI21_X1 port map( B1 => n168, B2 => n101, A => n119, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n108, ZN => n119);
   U60 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n118, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n101, ZN => n118);
   U62 : OAI21_X1 port map( B1 => n170, B2 => n101, A => n117, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => n101, ZN => n117);
   U64 : OAI21_X1 port map( B1 => n179, B2 => n108, A => n116, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n108, ZN => n116);
   U70 : CLKBUF_X1 port map( A => ld, Z => n101);
   U71 : CLKBUF_X1 port map( A => ld, Z => n102);
   U80 : CLKBUF_X1 port map( A => ld, Z => n108);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n179);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n178);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n177);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n176);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n175);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n174);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n173);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n172);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n171);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n170);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n169);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n168);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n167);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n166);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n165);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n164);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n163);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n162);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n161);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n160);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n159);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n158);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n157);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n156);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n155);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n154);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n153);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n152);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n151);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n150);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n149);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n148);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_10 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_10;

architecture SYN_behav of gen_reg_N32_10 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n100, n101, n102, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n161, B2 => n102, A => n137, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n100, A2 => data_in(23), ZN => n137);
   U4 : OAI21_X1 port map( B1 => n162, B2 => n102, A => n136, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n101, ZN => n136);
   U6 : OAI21_X1 port map( B1 => n163, B2 => n101, A => n135, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => n102, ZN => n135);
   U8 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n134, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => n100, ZN => n134);
   U10 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n133, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => n101, ZN => n133);
   U12 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n132, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => n102, ZN => n132);
   U14 : OAI21_X1 port map( B1 => n138, B2 => n101, A => n131, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => ld, ZN => n131);
   U16 : OAI21_X1 port map( B1 => n139, B2 => n100, A => n130, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n102, ZN => n130);
   U18 : OAI21_X1 port map( B1 => n140, B2 => n100, A => n129, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n129);
   U20 : OAI21_X1 port map( B1 => n167, B2 => n100, A => n128, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n101, ZN => n128);
   U22 : OAI21_X1 port map( B1 => n141, B2 => n100, A => n127, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n102, ZN => n127);
   U24 : OAI21_X1 port map( B1 => n142, B2 => n101, A => n126, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n102, ZN => n126);
   U26 : OAI21_X1 port map( B1 => n143, B2 => n100, A => n125, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n100, ZN => n125);
   U28 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n124, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => ld, ZN => n124);
   U30 : OAI21_X1 port map( B1 => n145, B2 => n101, A => n123, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n101, ZN => n123);
   U32 : OAI21_X1 port map( B1 => n146, B2 => n100, A => n122, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n101, ZN => n122);
   U34 : OAI21_X1 port map( B1 => n147, B2 => n100, A => n121, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n102, ZN => n121);
   U36 : OAI21_X1 port map( B1 => n148, B2 => n100, A => n120, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n101, ZN => n120);
   U38 : OAI21_X1 port map( B1 => n149, B2 => n100, A => n119, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n100, ZN => n119);
   U40 : OAI21_X1 port map( B1 => n150, B2 => n100, A => n118, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n100, ZN => n118);
   U42 : OAI21_X1 port map( B1 => n168, B2 => n100, A => n117, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => n101, ZN => n117);
   U44 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n116, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n100, ZN => n116);
   U46 : OAI21_X1 port map( B1 => n152, B2 => n100, A => n115, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => n102, ZN => n115);
   U48 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n114, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n102, ZN => n114);
   U50 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n113, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n102, ZN => n113);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n112, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n102, ZN => n112);
   U54 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n111, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n102, ZN => n111);
   U56 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n110, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n102, ZN => n110);
   U58 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n109, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n102, ZN => n109);
   U60 : OAI21_X1 port map( B1 => n159, B2 => n101, A => n108, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n102, ZN => n108);
   U62 : OAI21_X1 port map( B1 => n160, B2 => n102, A => n107, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => n102, ZN => n107);
   U64 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n106, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n100, ZN => n106);
   U72 : CLKBUF_X1 port map( A => ld, Z => n101);
   U73 : CLKBUF_X1 port map( A => ld, Z => n100);
   U74 : CLKBUF_X1 port map( A => ld, Z => n102);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n169);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n168);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n167);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n166);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n165);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n164);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n163);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n162);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n161);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n160);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n159);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n158);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n157);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n156);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n155);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n154);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n153);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n152);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n151);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n150);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n149);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n148);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n147);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n146);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n145);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n144);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n143);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n142);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n141);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n140);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n139);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n138);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_9 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_9;

architecture SYN_behav of gen_reg_N32_9 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n161, B2 => n97, A => n137, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n97, A2 => data_in(23), ZN => n137);
   U4 : OAI21_X1 port map( B1 => n162, B2 => n98, A => n136, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n136);
   U6 : OAI21_X1 port map( B1 => n163, B2 => ld, A => n135, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n135);
   U8 : OAI21_X1 port map( B1 => n164, B2 => ld, A => n134, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => n97, ZN => n134);
   U10 : OAI21_X1 port map( B1 => n165, B2 => ld, A => n133, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => ld, ZN => n133);
   U12 : OAI21_X1 port map( B1 => n166, B2 => n97, A => n132, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => n97, ZN => n132);
   U14 : OAI21_X1 port map( B1 => n138, B2 => ld, A => n131, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => n97, ZN => n131);
   U16 : OAI21_X1 port map( B1 => n139, B2 => n97, A => n130, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n98, ZN => n130);
   U18 : OAI21_X1 port map( B1 => n140, B2 => n98, A => n129, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n98, ZN => n129);
   U20 : OAI21_X1 port map( B1 => n167, B2 => n98, A => n128, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n128);
   U22 : OAI21_X1 port map( B1 => n141, B2 => ld, A => n127, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n98, ZN => n127);
   U24 : OAI21_X1 port map( B1 => n142, B2 => n98, A => n126, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n98, ZN => n126);
   U26 : OAI21_X1 port map( B1 => n143, B2 => ld, A => n125, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n98, ZN => n125);
   U28 : OAI21_X1 port map( B1 => n144, B2 => ld, A => n124, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n98, ZN => n124);
   U30 : OAI21_X1 port map( B1 => n145, B2 => n98, A => n123, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n98, ZN => n123);
   U32 : OAI21_X1 port map( B1 => n146, B2 => ld, A => n122, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n98, ZN => n122);
   U34 : OAI21_X1 port map( B1 => n147, B2 => ld, A => n121, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n98, ZN => n121);
   U36 : OAI21_X1 port map( B1 => n148, B2 => ld, A => n120, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n98, ZN => n120);
   U38 : OAI21_X1 port map( B1 => n149, B2 => ld, A => n119, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n98, ZN => n119);
   U40 : OAI21_X1 port map( B1 => n150, B2 => ld, A => n118, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n97, ZN => n118);
   U42 : OAI21_X1 port map( B1 => n168, B2 => ld, A => n117, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => n97, ZN => n117);
   U44 : OAI21_X1 port map( B1 => n151, B2 => ld, A => n116, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n97, ZN => n116);
   U46 : OAI21_X1 port map( B1 => n152, B2 => ld, A => n115, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => n97, ZN => n115);
   U48 : OAI21_X1 port map( B1 => n153, B2 => ld, A => n114, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n97, ZN => n114);
   U50 : OAI21_X1 port map( B1 => n154, B2 => ld, A => n113, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n97, ZN => n113);
   U52 : OAI21_X1 port map( B1 => n155, B2 => ld, A => n112, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n97, ZN => n112);
   U54 : OAI21_X1 port map( B1 => n156, B2 => ld, A => n111, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n97, ZN => n111);
   U56 : OAI21_X1 port map( B1 => n157, B2 => n97, A => n110, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n97, ZN => n110);
   U58 : OAI21_X1 port map( B1 => n158, B2 => ld, A => n109, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n97, ZN => n109);
   U60 : OAI21_X1 port map( B1 => n159, B2 => n98, A => n108, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n97, ZN => n108);
   U62 : OAI21_X1 port map( B1 => n160, B2 => n97, A => n107, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => n97, ZN => n107);
   U64 : OAI21_X1 port map( B1 => n169, B2 => n98, A => n106, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n98, ZN => n106);
   U69 : CLKBUF_X1 port map( A => ld, Z => n97);
   U70 : CLKBUF_X1 port map( A => ld, Z => n98);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n169);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n168);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n167);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n166);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n165);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n164);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n163);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n162);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n161);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n160);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n159);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n158);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n157);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n156);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n155);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n154);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n153);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n152);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n151);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n150);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n149);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n148);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n147);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n146);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n145);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n144);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n143);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n142);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n141);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n140);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n139);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n138);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_2 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_2;

architecture SYN_behav of gen_reg_N32_2 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n100, n102, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n161, B2 => n102, A => n137, ZN => n9);
   U3 : NAND2_X1 port map( A1 => ld, A2 => data_in(23), ZN => n137);
   U4 : OAI21_X1 port map( B1 => n162, B2 => n102, A => n136, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n102, ZN => n136);
   U6 : OAI21_X1 port map( B1 => n163, B2 => n102, A => n135, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => ld, ZN => n135);
   U8 : OAI21_X1 port map( B1 => n164, B2 => n100, A => n134, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => ld, ZN => n134);
   U10 : OAI21_X1 port map( B1 => n165, B2 => n102, A => n133, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => ld, ZN => n133);
   U12 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n132, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => ld, ZN => n132);
   U14 : OAI21_X1 port map( B1 => n138, B2 => n100, A => n131, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => ld, ZN => n131);
   U16 : OAI21_X1 port map( B1 => n139, B2 => n100, A => n130, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => ld, ZN => n130);
   U18 : OAI21_X1 port map( B1 => n140, B2 => n100, A => n129, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n100, ZN => n129);
   U20 : OAI21_X1 port map( B1 => n167, B2 => n100, A => n128, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => ld, ZN => n128);
   U22 : OAI21_X1 port map( B1 => n141, B2 => n100, A => n127, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => ld, ZN => n127);
   U24 : OAI21_X1 port map( B1 => n142, B2 => n100, A => n126, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => ld, ZN => n126);
   U26 : OAI21_X1 port map( B1 => n143, B2 => n100, A => n125, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => ld, ZN => n125);
   U28 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n124, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n102, ZN => n124);
   U30 : OAI21_X1 port map( B1 => n145, B2 => ld, A => n123, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n102, ZN => n123);
   U32 : OAI21_X1 port map( B1 => n146, B2 => n100, A => n122, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => ld, ZN => n122);
   U34 : OAI21_X1 port map( B1 => n147, B2 => n100, A => n121, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => ld, ZN => n121);
   U36 : OAI21_X1 port map( B1 => n148, B2 => n100, A => n120, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => ld, ZN => n120);
   U38 : OAI21_X1 port map( B1 => n149, B2 => n100, A => n119, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => ld, ZN => n119);
   U40 : OAI21_X1 port map( B1 => n150, B2 => n100, A => n118, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => ld, ZN => n118);
   U42 : OAI21_X1 port map( B1 => n168, B2 => n100, A => n117, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => n100, ZN => n117);
   U44 : OAI21_X1 port map( B1 => n151, B2 => n102, A => n116, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n100, ZN => n116);
   U46 : OAI21_X1 port map( B1 => n152, B2 => n100, A => n115, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => n102, ZN => n115);
   U48 : OAI21_X1 port map( B1 => n153, B2 => n100, A => n114, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n102, ZN => n114);
   U50 : OAI21_X1 port map( B1 => n154, B2 => n102, A => n113, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n102, ZN => n113);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n100, A => n112, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n102, ZN => n112);
   U54 : OAI21_X1 port map( B1 => n156, B2 => n102, A => n111, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n102, ZN => n111);
   U56 : OAI21_X1 port map( B1 => n157, B2 => n100, A => n110, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n102, ZN => n110);
   U58 : OAI21_X1 port map( B1 => n158, B2 => n102, A => n109, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n102, ZN => n109);
   U60 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n108, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n102, ZN => n108);
   U62 : OAI21_X1 port map( B1 => n160, B2 => n102, A => n107, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => n102, ZN => n107);
   U64 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n106, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n100, ZN => n106);
   U73 : CLKBUF_X1 port map( A => ld, Z => n100);
   U74 : CLKBUF_X1 port map( A => ld, Z => n102);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n169);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n168);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n167);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n166);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n165);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n164);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n163);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n162);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n161);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n160);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n159);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n158);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n157);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n156);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n155);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n154);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n153);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n152);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n151);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n150);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n149);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n148);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n147);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n146);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n145);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n144);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n143);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n142);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n141);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n140);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n139);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n138);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_1 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_1;

architecture SYN_behav of gen_reg_N32_1 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n100, n102, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n161, B2 => n102, A => n137, ZN => n9);
   U3 : NAND2_X1 port map( A1 => ld, A2 => data_in(23), ZN => n137);
   U4 : OAI21_X1 port map( B1 => n162, B2 => n102, A => n136, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n100, ZN => n136);
   U6 : OAI21_X1 port map( B1 => n163, B2 => n102, A => n135, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => ld, ZN => n135);
   U8 : OAI21_X1 port map( B1 => n164, B2 => n100, A => n134, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => ld, ZN => n134);
   U10 : OAI21_X1 port map( B1 => n165, B2 => n102, A => n133, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => ld, ZN => n133);
   U12 : OAI21_X1 port map( B1 => n166, B2 => n100, A => n132, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => ld, ZN => n132);
   U14 : OAI21_X1 port map( B1 => n138, B2 => n100, A => n131, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => ld, ZN => n131);
   U16 : OAI21_X1 port map( B1 => n139, B2 => n100, A => n130, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => ld, ZN => n130);
   U18 : OAI21_X1 port map( B1 => n140, B2 => n100, A => n129, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n102, ZN => n129);
   U20 : OAI21_X1 port map( B1 => n167, B2 => n100, A => n128, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => ld, ZN => n128);
   U22 : OAI21_X1 port map( B1 => n141, B2 => n100, A => n127, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => ld, ZN => n127);
   U24 : OAI21_X1 port map( B1 => n142, B2 => n100, A => n126, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => ld, ZN => n126);
   U26 : OAI21_X1 port map( B1 => n143, B2 => n100, A => n125, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => ld, ZN => n125);
   U28 : OAI21_X1 port map( B1 => n144, B2 => n102, A => n124, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => ld, ZN => n124);
   U30 : OAI21_X1 port map( B1 => n145, B2 => ld, A => n123, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => ld, ZN => n123);
   U32 : OAI21_X1 port map( B1 => n146, B2 => n100, A => n122, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => ld, ZN => n122);
   U34 : OAI21_X1 port map( B1 => n147, B2 => n100, A => n121, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => ld, ZN => n121);
   U36 : OAI21_X1 port map( B1 => n148, B2 => n100, A => n120, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => ld, ZN => n120);
   U38 : OAI21_X1 port map( B1 => n149, B2 => n100, A => n119, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => ld, ZN => n119);
   U40 : OAI21_X1 port map( B1 => n150, B2 => n100, A => n118, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => ld, ZN => n118);
   U42 : OAI21_X1 port map( B1 => n168, B2 => n100, A => n117, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => ld, ZN => n117);
   U44 : OAI21_X1 port map( B1 => n151, B2 => n102, A => n116, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => ld, ZN => n116);
   U46 : OAI21_X1 port map( B1 => n152, B2 => n100, A => n115, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => n102, ZN => n115);
   U48 : OAI21_X1 port map( B1 => n153, B2 => n100, A => n114, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n102, ZN => n114);
   U50 : OAI21_X1 port map( B1 => n154, B2 => n102, A => n113, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n102, ZN => n113);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n100, A => n112, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n102, ZN => n112);
   U54 : OAI21_X1 port map( B1 => n156, B2 => n102, A => n111, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n102, ZN => n111);
   U56 : OAI21_X1 port map( B1 => n157, B2 => n100, A => n110, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n102, ZN => n110);
   U58 : OAI21_X1 port map( B1 => n158, B2 => n102, A => n109, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n102, ZN => n109);
   U60 : OAI21_X1 port map( B1 => n159, B2 => n100, A => n108, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n102, ZN => n108);
   U62 : OAI21_X1 port map( B1 => n160, B2 => n102, A => n107, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => ld, ZN => n107);
   U64 : OAI21_X1 port map( B1 => n169, B2 => n102, A => n106, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => ld, ZN => n106);
   U73 : CLKBUF_X1 port map( A => ld, Z => n100);
   U74 : CLKBUF_X1 port map( A => ld, Z => n102);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n169);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n168);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n167);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n166);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n165);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n164);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n163);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n162);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n161);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n160);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n159);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n158);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n157);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n156);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n155);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n154);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n153);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n152);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n151);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n150);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n149);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n148);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n147);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n146);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n145);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n144);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n143);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n142);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n141);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n140);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n139);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n138);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N1_1 is

   port( clk, rst, ld, data_in : in std_logic;  data_out : out std_logic);

end gen_reg_N1_1;

architecture SYN_behav of gen_reg_N1_1 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n3, B2 => ld, A => n2, ZN => n1);
   U3 : NAND2_X1 port map( A1 => ld, A2 => data_in, ZN => n2);
   data_out_reg_0_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           data_out, QN => n3);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_add_0 is

   port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (29 downto 0);  CO : out std_logic);

end ALU_N32_DW01_add_0;

architecture SYN_cla of ALU_N32_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, n104, 
      n119, n121, n122, n129, n136, n140, n141, SUM_14_port, net82661, net82865
      , net82907, net82950, net82958, net83142, net83234, net83235, net83818, 
      net83800, net83773, net83772, net83767, net83859, net86251, net87686, 
      net87701, net87714, net88306, net88345, net88330, net88326, net96954, 
      net97018, net87770, net88944, net88378, net88367, net88354, net101217, 
      net101183, net101182, net101181, net110194, net110303, net110296, 
      net110294, net110284, net110237, net110236, net110331, net110344, 
      net110343, net110347, net99649, n135, n107, net118595, net118593, 
      net118590, net118557, net101208, net101201, net101193, net101191, 
      net101190, net101178, net101176, net118560, net118556, n105, net95105, 
      net88357, net88351, net118597, net118571, net101263, net101262, net101199
      , net101198, net101197, net101196, net101184, net101174, net96943, 
      net88964, net88963, net83837, net83836, net83835, net83834, net83832, 
      net83807, net83806, net83803, net83799, net118604, net118594, net83805, 
      net101195, net101188, net101186, net101156, net99637, net99634, net99631,
      net95069, net95068, net95054, net83879, net101310, net97049, net88307, 
      net83831, net83830, net83790, net83788, net83786, net101254, n75, n76, 
      n77, n82, n83, n85, n86, n87, n90, n91, n96, n97, n98, n99, n100, n101, 
      n102, n103, n106, n108, n109, n110, n112, n115, n116, n117, n120, n123, 
      n124, n128, n132, n133, n137, n138, n139, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168 : std_logic;

begin
   SUM <= ( SUM_29_port, SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_19_port, SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, 
      SUM_14_port, A(13), A(12), A(11), A(10), A(9), A(8), A(7), A(6), A(5), 
      A(4), A(3), A(2), A(1), A(0) );
   
   U16 : XOR2_X1 port map( A => B(14), B => net82661, Z => SUM_14_port);
   U56 : XNOR2_X1 port map( A => net83235, B => n122, ZN => SUM_20_port);
   U57 : NOR2_X1 port map( A1 => n119, A2 => net83790, ZN => n122);
   U58 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n121);
   U59 : NOR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n119);
   U65 : XNOR2_X1 port map( A => net82950, B => n129, ZN => SUM_18_port);
   U74 : XNOR2_X1 port map( A => n143, B => n136, ZN => SUM_16_port);
   U75 : NOR2_X1 port map( A1 => net82865, A2 => net95069, ZN => n136);
   U81 : XNOR2_X1 port map( A => n140, B => n141, ZN => SUM_15_port);
   U82 : NAND2_X1 port map( A1 => B(14), A2 => net82661, ZN => n141);
   U83 : AOI21_X1 port map( B1 => net87714, B2 => net82907, A => n137, ZN => 
                           n140);
   U76 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n135);
   U41 : NOR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n105);
   U40 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n107);
   U2 : OAI21_X1 port map( B1 => n75, B2 => n76, A => net88963, ZN => net83807)
                           ;
   U3 : NAND2_X1 port map( A1 => net101254, A2 => net83830, ZN => n75);
   U4 : INV_X1 port map( A => net96943, ZN => n76);
   U5 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n77);
   U15 : NAND2_X1 port map( A1 => net101184, A2 => net101190, ZN => n86);
   U18 : NAND2_X1 port map( A1 => n90, A2 => n154, ZN => n87);
   U20 : OR2_X1 port map( A1 => net88944, A2 => net110303, ZN => n90);
   U22 : NAND2_X1 port map( A1 => net83805, A2 => n148, ZN => n91);
   U23 : XNOR2_X1 port map( A => net83234, B => n146, ZN => SUM_21_port);
   U25 : XNOR2_X1 port map( A => n96, B => n150, ZN => SUM_29_port);
   U28 : AOI21_X1 port map( B1 => net101217, B2 => net87770, A => net101156, ZN
                           => net86251);
   U29 : INV_X1 port map( A => n105, ZN => net101217);
   U30 : INV_X1 port map( A => n107, ZN => net101156);
   U31 : NAND2_X1 port map( A1 => n132, A2 => net83859, ZN => net83800);
   U32 : AOI21_X1 port map( B1 => net101208, B2 => n144, A => n152, ZN => n96);
   U36 : NAND2_X1 port map( A1 => net101254, A2 => net96943, ZN => net118604);
   U37 : INV_X1 port map( A => A(19), ZN => net83788);
   U39 : AOI21_X1 port map( B1 => n168, B2 => net88357, A => n139, ZN => 
                           net88307);
   U43 : AOI21_X1 port map( B1 => net88351, B2 => net97049, A => n139, ZN => 
                           net88306);
   U44 : OR2_X1 port map( A1 => net83831, A2 => n121, ZN => net83830);
   U45 : INV_X1 port map( A => net83830, ZN => net88964);
   U46 : INV_X1 port map( A => A(21), ZN => net83831);
   U48 : CLKBUF_X1 port map( A => net110343, Z => net97049);
   U49 : AOI21_X1 port map( B1 => n138, B2 => net88357, A => n139, ZN => 
                           net83786);
   U51 : OAI21_X1 port map( B1 => net83235, B2 => n119, A => n121, ZN => 
                           net83234);
   U60 : NOR2_X1 port map( A1 => A(21), A2 => net83790, ZN => net83799);
   U63 : OR2_X1 port map( A1 => net95069, A2 => net99649, ZN => net95068);
   U66 : INV_X1 port map( A => n135, ZN => net95069);
   U67 : NAND2_X1 port map( A1 => net99631, A2 => B(14), ZN => net99634);
   U68 : NAND2_X1 port map( A1 => net99634, A2 => net95054, ZN => net101310);
   U69 : INV_X1 port map( A => net99637, ZN => net99631);
   U70 : NAND2_X1 port map( A1 => net99631, A2 => B(14), ZN => net110294);
   U71 : OAI21_X1 port map( B1 => A(15), B2 => B(15), A => A(14), ZN => 
                           net99637);
   U73 : AOI22_X1 port map( A1 => n161, A2 => net95054, B1 => net82865, B2 => 
                           n135, ZN => net110296);
   U77 : AOI22_X1 port map( A1 => net110294, A2 => net95054, B1 => net82865, B2
                           => n135, ZN => net95105);
   U78 : INV_X1 port map( A => net99649, ZN => net82865);
   U85 : CLKBUF_X1 port map( A => A(15), Z => net82907);
   U86 : NAND2_X1 port map( A1 => A(15), A2 => B(15), ZN => net83879);
   U87 : CLKBUF_X1 port map( A => B(15), Z => net87714);
   U88 : CLKBUF_X1 port map( A => A(14), Z => net82661);
   U94 : NOR2_X1 port map( A1 => B(25), A2 => net101156, ZN => n97);
   U96 : NAND2_X1 port map( A1 => n91, A2 => net87701, ZN => net87770);
   U99 : NAND2_X1 port map( A1 => net83807, A2 => net83806, ZN => net83805);
   U100 : NAND2_X1 port map( A1 => net101188, A2 => net101217, ZN => net101195)
                           ;
   U103 : NOR2_X1 port map( A1 => B(25), A2 => net101217, ZN => net101186);
   U104 : NAND2_X1 port map( A1 => n107, A2 => net101217, ZN => net96954);
   U106 : XNOR2_X1 port map( A => B(25), B => net101174, ZN => n104);
   U107 : NAND2_X1 port map( A1 => net101196, A2 => B(25), ZN => net101197);
   U109 : NAND2_X1 port map( A1 => net118560, A2 => net87686, ZN => net83773);
   U110 : NAND2_X1 port map( A1 => net118595, A2 => net118556, ZN => net118590)
                           ;
   U111 : NAND2_X1 port map( A1 => net118556, A2 => net118557, ZN => net87701);
   U113 : NAND2_X1 port map( A1 => n162, A2 => net83807, ZN => net87686);
   U114 : AOI21_X1 port map( B1 => n160, B2 => n162, A => net118590, ZN => 
                           net97018);
   U116 : NAND2_X1 port map( A1 => n105, A2 => n107, ZN => net118597);
   U117 : OR2_X1 port map( A1 => net88964, A2 => net83832, ZN => net88963);
   U119 : OR2_X1 port map( A1 => net83836, A2 => net83799, ZN => net83835);
   U120 : INV_X1 port map( A => B(21), ZN => net83836);
   U121 : NAND2_X1 port map( A1 => net83800, A2 => net83837, ZN => net83834);
   U124 : NAND2_X1 port map( A1 => net83832, A2 => net118604, ZN => net118594);
   U126 : OAI21_X1 port map( B1 => n98, B2 => n87, A => B(19), ZN => net96943);
   U130 : NAND2_X1 port map( A1 => n87, A2 => B(19), ZN => net110331);
   U132 : INV_X1 port map( A => net110296, ZN => net110284);
   U134 : NAND2_X1 port map( A1 => n77, A2 => A(17), ZN => net110194);
   U135 : NAND2_X1 port map( A1 => net101197, A2 => net101198, ZN => net101184)
                           ;
   U137 : INV_X1 port map( A => net101262, ZN => net101263);
   U138 : NAND2_X1 port map( A1 => net101199, A2 => A(25), ZN => net101262);
   U140 : AOI21_X1 port map( B1 => net118571, B2 => n162, A => n100, ZN => 
                           net101196);
   U141 : NAND2_X1 port map( A1 => n101, A2 => net118597, ZN => n100);
   U142 : NAND2_X1 port map( A1 => net118590, A2 => n107, ZN => n101);
   U143 : NOR2_X1 port map( A1 => net118593, A2 => net101156, ZN => net118571);
   U146 : NAND2_X1 port map( A1 => net110194, A2 => net88378, ZN => net88357);
   U148 : NAND2_X1 port map( A1 => net88354, A2 => net88944, ZN => n102);
   U150 : NAND2_X1 port map( A1 => net88378, A2 => net110194, ZN => net88351);
   U153 : INV_X1 port map( A => net88944, ZN => net88330);
   U154 : NAND2_X1 port map( A1 => n103, A2 => n106, ZN => net118560);
   U157 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => net118556);
   U160 : NAND2_X1 port map( A1 => n86, A2 => net101201, ZN => net101182);
   U161 : NAND2_X1 port map( A1 => net101176, A2 => net101178, ZN => net101190)
                           ;
   U162 : NAND2_X1 port map( A1 => net101190, A2 => net101201, ZN => net101183)
                           ;
   U169 : INV_X1 port map( A => A(27), ZN => net101193);
   U170 : NAND2_X1 port map( A1 => net101201, A2 => net101193, ZN => n112);
   U171 : INV_X1 port map( A => B(27), ZN => net101191);
   U172 : NAND2_X1 port map( A1 => net101201, A2 => net101191, ZN => n110);
   U174 : XNOR2_X1 port map( A => B(28), B => A(28), ZN => net83142);
   U175 : XNOR2_X1 port map( A => B(27), B => A(27), ZN => net101181);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => net101201);
   U179 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n115);
   U180 : NAND2_X1 port map( A1 => net83772, A2 => n115, ZN => net118557);
   U185 : NAND2_X1 port map( A1 => n117, A2 => n120, ZN => net110347);
   U186 : NAND2_X1 port map( A1 => net110343, A2 => net110344, ZN => n116);
   U188 : NAND2_X1 port map( A1 => n117, A2 => n120, ZN => net88367);
   U190 : NAND2_X1 port map( A1 => net88345, A2 => n123, ZN => net110236);
   U191 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => net110237);
   U192 : INV_X1 port map( A => A(18), ZN => n117);
   U193 : INV_X1 port map( A => B(18), ZN => n120);
   U195 : INV_X1 port map( A => A(17), ZN => net88345);
   U197 : XNOR2_X1 port map( A => net101182, B => net101181, ZN => SUM_27_port)
                           ;
   U198 : XNOR2_X1 port map( A => net101183, B => n124, ZN => SUM_26_port);
   U199 : NAND2_X1 port map( A1 => net101197, A2 => n164, ZN => n124);
   U201 : NAND2_X1 port map( A1 => B(17), A2 => net88367, ZN => net88378);
   U202 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => net88354);
   U203 : INV_X1 port map( A => net88354, ZN => net88326);
   U204 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => net88944);
   U206 : XNOR2_X1 port map( A => net97018, B => net96954, ZN => SUM_24_port);
   U212 : XNOR2_X1 port map( A => net87686, B => n128, ZN => SUM_22_port);
   U213 : OR2_X1 port map( A1 => net83767, A2 => n133, ZN => n128);
   U214 : NOR2_X1 port map( A1 => net88326, A2 => net110303, ZN => n129);
   U215 : AOI21_X1 port map( B1 => net110236, B2 => net110296, A => net88330, 
                           ZN => net82950);
   U217 : XNOR2_X1 port map( A => net110284, B => n151, ZN => SUM_17_port);
   U220 : INV_X1 port map( A => net83800, ZN => net83235);
   U221 : XNOR2_X1 port map( A => net82958, B => n147, ZN => SUM_23_port);
   U225 : XNOR2_X1 port map( A => net83818, B => n149, ZN => SUM_19_port);
   U227 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => net83772);
   U230 : INV_X1 port map( A => net88306, ZN => net83818);
   U232 : NAND2_X1 port map( A1 => net83773, A2 => net83772, ZN => net82958);
   U234 : NOR2_X1 port map( A1 => net87714, A2 => net82907, ZN => n137);
   U236 : XNOR2_X1 port map( A => net86251, B => n104, ZN => SUM_25_port);
   U6 : AND2_X1 port map( A1 => net83879, A2 => n135, ZN => net95054);
   U7 : OR2_X1 port map( A1 => net83786, A2 => net83788, ZN => net83859);
   U8 : OR2_X1 port map( A1 => net88307, A2 => net83788, ZN => net101254);
   U9 : AND2_X1 port map( A1 => net83834, A2 => net83835, ZN => n162);
   U10 : AOI22_X1 port map( A1 => net110294, A2 => net95054, B1 => net82865, B2
                           => n135, ZN => n138);
   U11 : AND2_X1 port map( A1 => n102, A2 => net110347, ZN => n139);
   U12 : OR2_X1 port map( A1 => A(27), A2 => B(27), ZN => n142);
   U13 : AND2_X1 port map( A1 => n161, A2 => net83879, ZN => n143);
   U14 : OR2_X1 port map( A1 => A(28), A2 => B(28), ZN => n144);
   U17 : AND2_X1 port map( A1 => net101195, A2 => n97, ZN => n145);
   U19 : XOR2_X1 port map( A => A(21), B => net83836, Z => n146);
   U21 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n147);
   U24 : AND2_X1 port map( A1 => net118560, A2 => net118556, ZN => n148);
   U26 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n149);
   U27 : XOR2_X1 port map( A => A(29), B => B(29), Z => n150);
   U33 : AND2_X1 port map( A1 => net110236, A2 => net110237, ZN => n151);
   U34 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n152);
   U35 : AND2_X1 port map( A1 => net83830, A2 => net87701, ZN => n153);
   U38 : AND2_X1 port map( A1 => net88354, A2 => net83788, ZN => n154);
   U42 : AND2_X1 port map( A1 => n112, A2 => n110, ZN => n155);
   U47 : NAND2_X1 port map( A1 => net83859, A2 => n159, ZN => n156);
   U50 : NAND2_X1 port map( A1 => n156, A2 => n157, ZN => net83806);
   U52 : OR2_X1 port map( A1 => n158, A2 => net83837, ZN => n157);
   U53 : INV_X1 port map( A => net83835, ZN => n158);
   U54 : AND2_X1 port map( A1 => n132, A2 => net83835, ZN => n159);
   U55 : NAND2_X1 port map( A1 => net118594, A2 => n153, ZN => net118593);
   U61 : AND3_X1 port map( A1 => net118594, A2 => net87701, A3 => net83830, ZN 
                           => n160);
   U62 : CLKBUF_X1 port map( A => net110294, Z => n161);
   U64 : XNOR2_X1 port map( A => n163, B => net83142, ZN => SUM_28_port);
   U72 : OR2_X1 port map( A1 => n83, A2 => n82, ZN => n163);
   U79 : OR2_X1 port map( A1 => n82, A2 => n83, ZN => net101208);
   U80 : AND2_X1 port map( A1 => n165, A2 => n166, ZN => n164);
   U84 : NAND2_X1 port map( A1 => net83805, A2 => n167, ZN => n165);
   U89 : AND2_X1 port map( A1 => n165, A2 => n166, ZN => net101198);
   U90 : OR2_X1 port map( A1 => net101262, A2 => n145, ZN => n166);
   U91 : AND2_X1 port map( A1 => n148, A2 => net101263, ZN => n167);
   U92 : AND2_X1 port map( A1 => net101310, A2 => net95068, ZN => n168);
   U93 : AND3_X1 port map( A1 => n77, A2 => B(19), A3 => net110236, ZN => 
                           net110344);
   U95 : AND2_X1 port map( A1 => net101190, A2 => n142, ZN => n85);
   U97 : AND2_X1 port map( A1 => net101310, A2 => net95068, ZN => net110343);
   U98 : INV_X1 port map( A => n119, ZN => net83803);
   U101 : INV_X1 port map( A => net87701, ZN => net101188);
   U102 : AND2_X1 port map( A1 => net83803, A2 => A(21), ZN => net83832);
   U105 : AND2_X1 port map( A1 => net95105, A2 => n99, ZN => n98);
   U108 : AND2_X1 port map( A1 => n77, A2 => net110236, ZN => n99);
   U112 : INV_X1 port map( A => B(22), ZN => n106);
   U115 : INV_X1 port map( A => A(22), ZN => n103);
   U118 : INV_X1 port map( A => B(23), ZN => n108);
   U122 : INV_X1 port map( A => A(23), ZN => n109);
   U123 : AND2_X1 port map( A1 => n142, A2 => n155, ZN => n83);
   U125 : AND2_X1 port map( A1 => net101184, A2 => n85, ZN => n82);
   U127 : INV_X1 port map( A => net118560, ZN => net83767);
   U128 : AND2_X1 port map( A1 => n117, A2 => n120, ZN => net110303);
   U129 : OR2_X1 port map( A1 => A(16), A2 => B(16), ZN => net99649);
   U131 : INV_X1 port map( A => B(17), ZN => n123);
   U133 : INV_X1 port map( A => n121, ZN => net83790);
   U136 : AND2_X1 port map( A1 => net83803, A2 => B(21), ZN => net83837);
   U139 : AND2_X1 port map( A1 => n116, A2 => net110331, ZN => n132);
   U144 : NAND3_X1 port map( A1 => n107, A2 => net101186, A3 => net101195, ZN 
                           => net101199);
   U145 : NAND3_X1 port map( A1 => n115, A2 => net83767, A3 => net83772, ZN => 
                           net118595);
   U147 : INV_X1 port map( A => A(25), ZN => net101174);
   U149 : INV_X1 port map( A => B(26), ZN => net101178);
   U151 : INV_X1 port map( A => A(26), ZN => net101176);
   U152 : INV_X1 port map( A => net83772, ZN => n133);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW02_mult_0 is

   port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (31 downto 0));

end ALU_N32_DW02_mult_0;

architecture SYN_csa of ALU_N32_DW02_mult_0 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ALU_N32_DW01_add_0
      port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (29 downto 0);  CO : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal ab_15_15_port, ab_15_14_port, ab_15_13_port, ab_15_12_port, 
      ab_15_11_port, ab_15_10_port, ab_15_9_port, ab_15_8_port, ab_15_7_port, 
      ab_15_6_port, ab_15_5_port, ab_15_4_port, ab_15_3_port, ab_15_2_port, 
      ab_15_1_port, ab_15_0_port, ab_14_15_port, ab_14_14_port, ab_14_13_port, 
      ab_14_12_port, ab_14_11_port, ab_14_10_port, ab_14_9_port, ab_14_8_port, 
      ab_14_7_port, ab_14_6_port, ab_14_5_port, ab_14_4_port, ab_14_3_port, 
      ab_14_2_port, ab_14_1_port, ab_14_0_port, ab_13_15_port, ab_13_14_port, 
      ab_13_13_port, ab_13_12_port, ab_13_11_port, ab_13_10_port, ab_13_9_port,
      ab_13_8_port, ab_13_7_port, ab_13_6_port, ab_13_5_port, ab_13_4_port, 
      ab_13_3_port, ab_13_2_port, ab_13_1_port, ab_13_0_port, ab_12_15_port, 
      ab_12_14_port, ab_12_13_port, ab_12_12_port, ab_12_11_port, ab_12_10_port
      , ab_12_9_port, ab_12_8_port, ab_12_7_port, ab_12_6_port, ab_12_5_port, 
      ab_12_4_port, ab_12_3_port, ab_12_2_port, ab_12_1_port, ab_12_0_port, 
      ab_11_15_port, ab_11_14_port, ab_11_13_port, ab_11_12_port, ab_11_11_port
      , ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port, ab_11_6_port, 
      ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, ab_11_1_port, 
      ab_11_0_port, ab_10_15_port, ab_10_14_port, ab_10_13_port, ab_10_12_port,
      ab_10_11_port, ab_10_10_port, ab_10_9_port, ab_10_8_port, ab_10_7_port, 
      ab_10_6_port, ab_10_5_port, ab_10_4_port, ab_10_3_port, ab_10_2_port, 
      ab_10_1_port, ab_10_0_port, ab_9_15_port, ab_9_14_port, ab_9_13_port, 
      ab_9_12_port, ab_9_11_port, ab_9_10_port, ab_9_9_port, ab_9_8_port, 
      ab_9_6_port, ab_9_5_port, ab_9_4_port, ab_9_3_port, ab_9_2_port, 
      ab_9_1_port, ab_9_0_port, ab_8_15_port, ab_8_14_port, ab_8_13_port, 
      ab_8_12_port, ab_8_11_port, ab_8_10_port, ab_8_9_port, ab_8_8_port, 
      ab_8_7_port, ab_8_6_port, ab_8_5_port, ab_8_4_port, ab_8_3_port, 
      ab_8_2_port, ab_8_1_port, ab_8_0_port, ab_7_15_port, ab_7_14_port, 
      ab_7_13_port, ab_7_12_port, ab_7_11_port, ab_7_10_port, ab_7_9_port, 
      ab_7_8_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_15_port, 
      ab_6_14_port, ab_6_13_port, ab_6_12_port, ab_6_11_port, ab_6_10_port, 
      ab_6_9_port, ab_6_8_port, ab_6_7_port, ab_6_6_port, ab_6_5_port, 
      ab_6_4_port, ab_6_3_port, ab_6_2_port, ab_6_1_port, ab_6_0_port, 
      ab_5_15_port, ab_5_14_port, ab_5_13_port, ab_5_12_port, ab_5_11_port, 
      ab_5_9_port, ab_5_8_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_15_port, ab_4_14_port, ab_4_13_port, ab_4_12_port, ab_4_11_port, 
      ab_4_10_port, ab_4_9_port, ab_4_8_port, ab_4_7_port, ab_4_6_port, 
      ab_4_5_port, ab_4_4_port, ab_4_3_port, ab_4_2_port, ab_4_1_port, 
      ab_4_0_port, ab_3_15_port, ab_3_14_port, ab_3_13_port, ab_3_12_port, 
      ab_3_10_port, ab_3_9_port, ab_3_8_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_15_port, ab_2_14_port, ab_2_13_port, ab_2_11_port, 
      ab_2_10_port, ab_2_9_port, ab_2_8_port, ab_2_7_port, ab_2_6_port, 
      ab_2_5_port, ab_2_4_port, ab_2_3_port, ab_2_2_port, ab_2_1_port, 
      ab_2_0_port, ab_1_15_port, ab_1_11_port, ab_1_10_port, ab_1_9_port, 
      ab_1_7_port, ab_1_6_port, ab_1_5_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_12_port, ab_0_11_port, ab_0_10_port, 
      ab_0_9_port, ab_0_8_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_15_15_port, 
      CARRYB_15_14_port, CARRYB_15_13_port, CARRYB_15_12_port, 
      CARRYB_15_11_port, CARRYB_15_10_port, CARRYB_15_9_port, CARRYB_15_8_port,
      CARRYB_15_7_port, CARRYB_15_6_port, CARRYB_15_5_port, CARRYB_15_4_port, 
      CARRYB_15_3_port, CARRYB_15_2_port, CARRYB_15_0_port, CARRYB_14_14_port, 
      CARRYB_14_13_port, CARRYB_14_12_port, CARRYB_14_11_port, 
      CARRYB_14_10_port, CARRYB_14_9_port, CARRYB_14_8_port, CARRYB_14_7_port, 
      CARRYB_14_6_port, CARRYB_14_5_port, CARRYB_14_4_port, CARRYB_14_3_port, 
      CARRYB_14_1_port, CARRYB_14_0_port, CARRYB_13_14_port, CARRYB_13_13_port,
      CARRYB_13_12_port, CARRYB_13_11_port, CARRYB_13_10_port, CARRYB_13_9_port
      , CARRYB_13_8_port, CARRYB_13_7_port, CARRYB_13_6_port, CARRYB_13_5_port,
      CARRYB_13_4_port, CARRYB_13_2_port, CARRYB_13_1_port, CARRYB_13_0_port, 
      CARRYB_12_14_port, CARRYB_12_13_port, CARRYB_12_12_port, 
      CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port, CARRYB_12_8_port,
      CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port, CARRYB_12_2_port, 
      CARRYB_12_1_port, CARRYB_12_0_port, CARRYB_11_14_port, CARRYB_11_13_port,
      CARRYB_11_12_port, CARRYB_11_11_port, CARRYB_11_10_port, CARRYB_11_9_port
      , CARRYB_11_8_port, CARRYB_11_7_port, CARRYB_11_6_port, CARRYB_11_2_port,
      CARRYB_11_1_port, CARRYB_11_0_port, CARRYB_10_14_port, CARRYB_10_13_port,
      CARRYB_10_12_port, CARRYB_10_11_port, CARRYB_10_10_port, CARRYB_10_9_port
      , CARRYB_10_8_port, CARRYB_10_7_port, CARRYB_10_3_port, CARRYB_10_2_port,
      CARRYB_10_1_port, CARRYB_10_0_port, CARRYB_9_14_port, CARRYB_9_13_port, 
      CARRYB_9_12_port, CARRYB_9_11_port, CARRYB_9_10_port, CARRYB_9_9_port, 
      CARRYB_9_8_port, CARRYB_9_4_port, CARRYB_9_3_port, CARRYB_9_2_port, 
      CARRYB_9_1_port, CARRYB_9_0_port, CARRYB_8_14_port, CARRYB_8_13_port, 
      CARRYB_8_12_port, CARRYB_8_11_port, CARRYB_8_10_port, CARRYB_8_9_port, 
      CARRYB_8_8_port, CARRYB_8_5_port, CARRYB_8_4_port, CARRYB_8_3_port, 
      CARRYB_8_2_port, CARRYB_8_1_port, CARRYB_8_0_port, CARRYB_7_14_port, 
      CARRYB_7_13_port, CARRYB_7_12_port, CARRYB_7_11_port, CARRYB_7_10_port, 
      CARRYB_7_9_port, CARRYB_7_6_port, CARRYB_7_5_port, CARRYB_7_4_port, 
      CARRYB_7_3_port, CARRYB_7_2_port, CARRYB_7_1_port, CARRYB_7_0_port, 
      CARRYB_6_14_port, CARRYB_6_13_port, CARRYB_6_12_port, CARRYB_6_11_port, 
      CARRYB_6_10_port, CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_14_port, CARRYB_5_13_port, CARRYB_5_12_port, 
      CARRYB_5_11_port, CARRYB_5_8_port, CARRYB_5_7_port, CARRYB_5_6_port, 
      CARRYB_5_5_port, CARRYB_5_4_port, CARRYB_5_3_port, CARRYB_5_2_port, 
      CARRYB_5_1_port, CARRYB_5_0_port, CARRYB_4_14_port, CARRYB_4_13_port, 
      CARRYB_4_12_port, CARRYB_4_11_port, CARRYB_4_9_port, CARRYB_4_8_port, 
      CARRYB_4_7_port, CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, 
      CARRYB_4_3_port, CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, 
      CARRYB_3_14_port, CARRYB_3_13_port, CARRYB_3_12_port, CARRYB_3_10_port, 
      CARRYB_3_9_port, CARRYB_3_8_port, CARRYB_3_7_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_14_port, CARRYB_2_13_port, 
      CARRYB_2_11_port, CARRYB_2_10_port, CARRYB_2_9_port, CARRYB_2_8_port, 
      CARRYB_2_7_port, CARRYB_2_6_port, CARRYB_2_5_port, CARRYB_2_4_port, 
      CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, CARRYB_2_0_port, 
      SUMB_15_15_port, SUMB_15_14_port, SUMB_15_13_port, SUMB_15_12_port, 
      SUMB_15_11_port, SUMB_15_10_port, SUMB_15_9_port, SUMB_15_8_port, 
      SUMB_15_7_port, SUMB_15_6_port, SUMB_15_5_port, SUMB_15_4_port, 
      SUMB_15_3_port, SUMB_15_2_port, SUMB_15_0_port, SUMB_14_14_port, 
      SUMB_14_13_port, SUMB_14_12_port, SUMB_14_11_port, SUMB_14_10_port, 
      SUMB_14_9_port, SUMB_14_8_port, SUMB_14_7_port, SUMB_14_6_port, 
      SUMB_14_5_port, SUMB_14_4_port, SUMB_14_3_port, SUMB_14_1_port, 
      SUMB_13_14_port, SUMB_13_13_port, SUMB_13_12_port, SUMB_13_11_port, 
      SUMB_13_10_port, SUMB_13_9_port, SUMB_13_8_port, SUMB_13_7_port, 
      SUMB_13_6_port, SUMB_13_5_port, SUMB_13_2_port, SUMB_13_1_port, 
      SUMB_12_14_port, SUMB_12_13_port, SUMB_12_12_port, SUMB_12_11_port, 
      SUMB_12_10_port, SUMB_12_9_port, SUMB_12_8_port, SUMB_12_7_port, 
      SUMB_12_6_port, SUMB_12_5_port, SUMB_12_2_port, SUMB_12_1_port, 
      SUMB_11_14_port, SUMB_11_13_port, SUMB_11_12_port, SUMB_11_11_port, 
      SUMB_11_10_port, SUMB_11_9_port, SUMB_11_8_port, SUMB_11_7_port, 
      SUMB_11_6_port, SUMB_11_2_port, SUMB_11_1_port, SUMB_10_14_port, 
      SUMB_10_13_port, SUMB_10_12_port, SUMB_10_11_port, SUMB_10_10_port, 
      SUMB_10_9_port, SUMB_10_8_port, SUMB_10_7_port, SUMB_10_3_port, 
      SUMB_10_2_port, SUMB_10_1_port, SUMB_9_14_port, SUMB_9_13_port, 
      SUMB_9_12_port, SUMB_9_11_port, SUMB_9_10_port, SUMB_9_9_port, 
      SUMB_9_8_port, SUMB_9_4_port, SUMB_9_3_port, SUMB_9_2_port, SUMB_9_1_port
      , SUMB_8_14_port, SUMB_8_13_port, SUMB_8_12_port, SUMB_8_11_port, 
      SUMB_8_10_port, SUMB_8_9_port, SUMB_8_5_port, SUMB_8_4_port, 
      SUMB_8_3_port, SUMB_8_2_port, SUMB_8_1_port, SUMB_7_14_port, 
      SUMB_7_13_port, SUMB_7_12_port, SUMB_7_11_port, SUMB_7_10_port, 
      SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, SUMB_7_3_port, SUMB_7_2_port
      , SUMB_7_1_port, SUMB_6_14_port, SUMB_6_13_port, SUMB_6_12_port, 
      SUMB_6_11_port, SUMB_6_10_port, SUMB_6_7_port, SUMB_6_6_port, 
      SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, SUMB_6_1_port
      , SUMB_5_14_port, SUMB_5_13_port, SUMB_5_12_port, SUMB_5_11_port, 
      SUMB_5_8_port, SUMB_5_7_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port
      , SUMB_5_3_port, SUMB_5_2_port, SUMB_5_1_port, SUMB_4_14_port, 
      SUMB_4_13_port, SUMB_4_12_port, SUMB_4_9_port, SUMB_4_8_port, 
      SUMB_4_7_port, SUMB_4_6_port, SUMB_4_5_port, SUMB_4_4_port, SUMB_4_3_port
      , SUMB_4_2_port, SUMB_4_1_port, SUMB_3_14_port, SUMB_3_13_port, 
      SUMB_3_12_port, SUMB_3_10_port, SUMB_3_9_port, SUMB_3_8_port, 
      SUMB_3_7_port, SUMB_3_6_port, SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port
      , SUMB_3_2_port, SUMB_3_1_port, SUMB_2_14_port, SUMB_2_13_port, 
      SUMB_2_11_port, SUMB_2_10_port, SUMB_2_9_port, SUMB_2_8_port, 
      SUMB_2_7_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, QA, QB, ZA, A1_13_port, A1_12_port, 
      A1_11_port, A1_10_port, A1_9_port, A1_8_port, A1_7_port, A1_6_port, 
      A1_5_port, A1_4_port, A1_3_port, A1_2_port, A1_1_port, A1_0_port, 
      A2_14_port, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n34, 
      n35, n36, n37, n38, n39, n40, n41, n49, n50, n51, n52, n53, n54, n62, n63
      , n98, n99, n61, n60, n59, n58, n57, n56, n55, n48, n47, n46, n45, n44, 
      n43, n42, n32, n100, n101, net74664, net74665, net74669, net74673, 
      net74680, net74690, net74691, net74693, net74694, net76791, net77069, 
      net77076, net77075, net82309, net82387, net82385, net82414, net82441, 
      net82475, net82535, net82597, net82595, net82608, net82622, net82635, 
      net82633, net82653, net82681, net82679, net82724, net82767, net82778, 
      net82876, net82942, net82976, net82975, net82980, net82987, net83062, 
      net83064, net83102, net83939, net83937, net83936, net86250, net86248, 
      net86247, net86245, net86243, net88957, net88956, net88955, net92268, 
      net92266, net95080, net96980, net97008, net118627, net118631, net118629, 
      net97026, SUMB_15_1_port, CARRYB_15_1_port, net82396, ab_5_10_port, 
      SUMB_4_11_port, SUMB_12_3_port, CARRYB_9_6_port, CARRYB_8_7_port, 
      CARRYB_7_8_port, CARRYB_6_9_port, CARRYB_5_10_port, CARRYB_12_3_port, 
      CARRYB_11_4_port, CARRYB_10_5_port, SUMB_11_4_port, SUMB_11_3_port, 
      CARRYB_11_3_port, net82986, ab_0_13_port, SUMB_14_2_port, 
      CARRYB_14_2_port, net82505, net74687, ab_9_7_port, SUMB_9_7_port, 
      SUMB_8_8_port, SUMB_7_9_port, SUMB_13_3_port, SUMB_12_4_port, 
      SUMB_11_5_port, SUMB_10_6_port, CARRYB_9_7_port, CARRYB_13_3_port, 
      CARRYB_12_4_port, CARRYB_11_5_port, CARRYB_10_6_port, SUMB_10_5_port, 
      SUMB_10_4_port, CARRYB_10_4_port, SUMB_9_6_port, SUMB_9_5_port, 
      CARRYB_9_5_port, SUMB_8_7_port, SUMB_8_6_port, CARRYB_8_6_port, 
      SUMB_7_8_port, SUMB_7_7_port, CARRYB_7_7_port, SUMB_6_9_port, 
      SUMB_6_8_port, CARRYB_6_8_port, SUMB_5_9_port, SUMB_5_10_port, 
      CARRYB_5_9_port, SUMB_4_10_port, CARRYB_4_10_port, net82716, net82651, 
      net74692, net74666, n26, n11, ab_3_11_port, ab_2_12_port, ab_1_12_port, 
      SUMB_3_11_port, SUMB_2_12_port, CARRYB_3_11_port, CARRYB_2_12_port, 
      net83044, net82534, n102, n105, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n161, n162, n163, n166, n167, n168, 
      n170, n171, n172, n173, n174, n175, n176, n177, n181, n184, n185, n186, 
      n187, n189, n192, n194, n197, n198, n199, n200, n201, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n238, n239, n240, n241, n242, n243, n245, n248, n265, 
      n266, n267, n272, n274, n275, n276, n278, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n_1020 : 
      std_logic;

begin
   
   S4_6 : FA_X1 port map( A => ab_15_6_port, B => CARRYB_14_6_port, CI => 
                           SUMB_14_7_port, CO => CARRYB_15_6_port, S => 
                           SUMB_15_6_port);
   S4_7 : FA_X1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, CI => 
                           SUMB_14_8_port, CO => CARRYB_15_7_port, S => 
                           SUMB_15_7_port);
   S4_8 : FA_X1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, CI => 
                           SUMB_14_9_port, CO => CARRYB_15_8_port, S => 
                           SUMB_15_8_port);
   S4_9 : FA_X1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, CI => 
                           SUMB_14_10_port, CO => CARRYB_15_9_port, S => 
                           SUMB_15_9_port);
   S4_10 : FA_X1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, CI => 
                           SUMB_14_11_port, CO => CARRYB_15_10_port, S => 
                           SUMB_15_10_port);
   S4_11 : FA_X1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, CI => 
                           SUMB_14_12_port, CO => CARRYB_15_11_port, S => 
                           SUMB_15_11_port);
   S4_12 : FA_X1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, CI => 
                           SUMB_14_13_port, CO => CARRYB_15_12_port, S => 
                           SUMB_15_12_port);
   S4_13 : FA_X1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, CI => 
                           SUMB_14_14_port, CO => CARRYB_15_13_port, S => 
                           SUMB_15_13_port);
   S5_14 : FA_X1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, CI => 
                           ab_14_15_port, CO => CARRYB_15_14_port, S => 
                           SUMB_15_14_port);
   S14_15 : FA_X1 port map( A => QA, B => QB, CI => ab_15_15_port, CO => 
                           CARRYB_15_15_port, S => SUMB_15_15_port);
   S2_14_1 : FA_X1 port map( A => CARRYB_13_1_port, B => ab_14_1_port, CI => 
                           SUMB_13_2_port, CO => CARRYB_14_1_port, S => 
                           SUMB_14_1_port);
   S2_14_4 : FA_X1 port map( A => ab_14_4_port, B => CARRYB_13_4_port, CI => 
                           SUMB_13_5_port, CO => CARRYB_14_4_port, S => 
                           SUMB_14_4_port);
   S2_14_7 : FA_X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, CI => 
                           SUMB_13_8_port, CO => CARRYB_14_7_port, S => 
                           SUMB_14_7_port);
   S2_14_8 : FA_X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, CI => 
                           SUMB_13_9_port, CO => CARRYB_14_8_port, S => 
                           SUMB_14_8_port);
   S2_14_9 : FA_X1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, CI => 
                           SUMB_13_10_port, CO => CARRYB_14_9_port, S => 
                           SUMB_14_9_port);
   S2_14_10 : FA_X1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, CI =>
                           SUMB_13_11_port, CO => CARRYB_14_10_port, S => 
                           SUMB_14_10_port);
   S2_14_11 : FA_X1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, CI =>
                           SUMB_13_12_port, CO => CARRYB_14_11_port, S => 
                           SUMB_14_11_port);
   S2_14_12 : FA_X1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, CI =>
                           SUMB_13_13_port, CO => CARRYB_14_12_port, S => 
                           SUMB_14_12_port);
   S2_14_13 : FA_X1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, CI =>
                           SUMB_13_14_port, CO => CARRYB_14_13_port, S => 
                           SUMB_14_13_port);
   S3_14_14 : FA_X1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, CI =>
                           ab_13_15_port, CO => CARRYB_14_14_port, S => 
                           SUMB_14_14_port);
   S1_13_0 : FA_X1 port map( A => CARRYB_12_0_port, B => ab_13_0_port, CI => 
                           SUMB_12_1_port, CO => CARRYB_13_0_port, S => 
                           A1_11_port);
   S2_13_1 : FA_X1 port map( A => CARRYB_12_1_port, B => ab_13_1_port, CI => 
                           SUMB_12_2_port, CO => CARRYB_13_1_port, S => 
                           SUMB_13_1_port);
   S2_13_5 : FA_X1 port map( A => ab_13_5_port, B => CARRYB_12_5_port, CI => 
                           SUMB_12_6_port, CO => CARRYB_13_5_port, S => 
                           SUMB_13_5_port);
   S2_13_7 : FA_X1 port map( A => CARRYB_12_7_port, B => ab_13_7_port, CI => 
                           SUMB_12_8_port, CO => CARRYB_13_7_port, S => 
                           SUMB_13_7_port);
   S2_13_8 : FA_X1 port map( A => ab_13_8_port, B => CARRYB_12_8_port, CI => 
                           SUMB_12_9_port, CO => CARRYB_13_8_port, S => 
                           SUMB_13_8_port);
   S2_13_9 : FA_X1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, CI => 
                           SUMB_12_10_port, CO => CARRYB_13_9_port, S => 
                           SUMB_13_9_port);
   S2_13_10 : FA_X1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, CI =>
                           SUMB_12_11_port, CO => CARRYB_13_10_port, S => 
                           SUMB_13_10_port);
   S2_13_11 : FA_X1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, CI =>
                           SUMB_12_12_port, CO => CARRYB_13_11_port, S => 
                           SUMB_13_11_port);
   S2_13_12 : FA_X1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, CI =>
                           SUMB_12_13_port, CO => CARRYB_13_12_port, S => 
                           SUMB_13_12_port);
   S2_13_13 : FA_X1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, CI =>
                           SUMB_12_14_port, CO => CARRYB_13_13_port, S => 
                           SUMB_13_13_port);
   S3_13_14 : FA_X1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, CI =>
                           ab_12_15_port, CO => CARRYB_13_14_port, S => 
                           SUMB_13_14_port);
   S1_12_0 : FA_X1 port map( A => CARRYB_11_0_port, B => ab_12_0_port, CI => 
                           SUMB_11_1_port, CO => CARRYB_12_0_port, S => 
                           A1_10_port);
   S2_12_1 : FA_X1 port map( A => CARRYB_11_1_port, B => ab_12_1_port, CI => 
                           SUMB_11_2_port, CO => CARRYB_12_1_port, S => 
                           SUMB_12_1_port);
   S2_12_8 : FA_X1 port map( A => CARRYB_11_8_port, B => ab_12_8_port, CI => 
                           SUMB_11_9_port, CO => CARRYB_12_8_port, S => 
                           SUMB_12_8_port);
   S2_12_9 : FA_X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, CI => 
                           SUMB_11_10_port, CO => CARRYB_12_9_port, S => 
                           SUMB_12_9_port);
   S2_12_10 : FA_X1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, CI =>
                           SUMB_11_11_port, CO => CARRYB_12_10_port, S => 
                           SUMB_12_10_port);
   S2_12_11 : FA_X1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, CI =>
                           SUMB_11_12_port, CO => CARRYB_12_11_port, S => 
                           SUMB_12_11_port);
   S2_12_12 : FA_X1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, CI =>
                           SUMB_11_13_port, CO => CARRYB_12_12_port, S => 
                           SUMB_12_12_port);
   S2_12_13 : FA_X1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, CI =>
                           SUMB_11_14_port, CO => CARRYB_12_13_port, S => 
                           SUMB_12_13_port);
   S3_12_14 : FA_X1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, CI =>
                           ab_11_15_port, CO => CARRYB_12_14_port, S => 
                           SUMB_12_14_port);
   S1_11_0 : FA_X1 port map( A => ab_11_0_port, B => CARRYB_10_0_port, CI => 
                           SUMB_10_1_port, CO => CARRYB_11_0_port, S => 
                           A1_9_port);
   S2_11_1 : FA_X1 port map( A => CARRYB_10_1_port, B => ab_11_1_port, CI => 
                           SUMB_10_2_port, CO => CARRYB_11_1_port, S => 
                           SUMB_11_1_port);
   S2_11_2 : FA_X1 port map( A => CARRYB_10_2_port, B => ab_11_2_port, CI => 
                           SUMB_10_3_port, CO => CARRYB_11_2_port, S => 
                           SUMB_11_2_port);
   S2_11_8 : FA_X1 port map( A => ab_11_8_port, B => CARRYB_10_8_port, CI => 
                           SUMB_10_9_port, CO => CARRYB_11_8_port, S => 
                           SUMB_11_8_port);
   S2_11_9 : FA_X1 port map( A => CARRYB_10_9_port, B => ab_11_9_port, CI => 
                           SUMB_10_10_port, CO => CARRYB_11_9_port, S => 
                           SUMB_11_9_port);
   S2_11_10 : FA_X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, CI =>
                           SUMB_10_11_port, CO => CARRYB_11_10_port, S => 
                           SUMB_11_10_port);
   S2_11_11 : FA_X1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, CI =>
                           SUMB_10_12_port, CO => CARRYB_11_11_port, S => 
                           SUMB_11_11_port);
   S2_11_12 : FA_X1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, CI =>
                           SUMB_10_13_port, CO => CARRYB_11_12_port, S => 
                           SUMB_11_12_port);
   S2_11_13 : FA_X1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, CI =>
                           SUMB_10_14_port, CO => CARRYB_11_13_port, S => 
                           SUMB_11_13_port);
   S3_11_14 : FA_X1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, CI =>
                           ab_10_15_port, CO => CARRYB_11_14_port, S => 
                           SUMB_11_14_port);
   S1_10_0 : FA_X1 port map( A => ab_10_0_port, B => CARRYB_9_0_port, CI => 
                           SUMB_9_1_port, CO => CARRYB_10_0_port, S => 
                           A1_8_port);
   S2_10_1 : FA_X1 port map( A => CARRYB_9_1_port, B => ab_10_1_port, CI => 
                           SUMB_9_2_port, CO => CARRYB_10_1_port, S => 
                           SUMB_10_1_port);
   S2_10_2 : FA_X1 port map( A => CARRYB_9_2_port, B => ab_10_2_port, CI => 
                           SUMB_9_3_port, CO => CARRYB_10_2_port, S => 
                           SUMB_10_2_port);
   S2_10_3 : FA_X1 port map( A => CARRYB_9_3_port, B => ab_10_3_port, CI => 
                           SUMB_9_4_port, CO => CARRYB_10_3_port, S => 
                           SUMB_10_3_port);
   S2_10_9 : FA_X1 port map( A => ab_10_9_port, B => CARRYB_9_9_port, CI => 
                           SUMB_9_10_port, CO => CARRYB_10_9_port, S => 
                           SUMB_10_9_port);
   S2_10_10 : FA_X1 port map( A => CARRYB_9_10_port, B => ab_10_10_port, CI => 
                           SUMB_9_11_port, CO => CARRYB_10_10_port, S => 
                           SUMB_10_10_port);
   S2_10_11 : FA_X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, CI => 
                           SUMB_9_12_port, CO => CARRYB_10_11_port, S => 
                           SUMB_10_11_port);
   S2_10_12 : FA_X1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, CI => 
                           SUMB_9_13_port, CO => CARRYB_10_12_port, S => 
                           SUMB_10_12_port);
   S2_10_13 : FA_X1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, CI => 
                           SUMB_9_14_port, CO => CARRYB_10_13_port, S => 
                           SUMB_10_13_port);
   S3_10_14 : FA_X1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, CI => 
                           ab_9_15_port, CO => CARRYB_10_14_port, S => 
                           SUMB_10_14_port);
   S1_9_0 : FA_X1 port map( A => ab_9_0_port, B => CARRYB_8_0_port, CI => 
                           SUMB_8_1_port, CO => CARRYB_9_0_port, S => A1_7_port
                           );
   S2_9_1 : FA_X1 port map( A => CARRYB_8_1_port, B => ab_9_1_port, CI => 
                           SUMB_8_2_port, CO => CARRYB_9_1_port, S => 
                           SUMB_9_1_port);
   S2_9_2 : FA_X1 port map( A => ab_9_2_port, B => CARRYB_8_2_port, CI => 
                           SUMB_8_3_port, CO => CARRYB_9_2_port, S => 
                           SUMB_9_2_port);
   S2_9_3 : FA_X1 port map( A => CARRYB_8_3_port, B => ab_9_3_port, CI => 
                           SUMB_8_4_port, CO => CARRYB_9_3_port, S => 
                           SUMB_9_3_port);
   S2_9_4 : FA_X1 port map( A => CARRYB_8_4_port, B => ab_9_4_port, CI => 
                           SUMB_8_5_port, CO => CARRYB_9_4_port, S => 
                           SUMB_9_4_port);
   S2_9_8 : FA_X1 port map( A => ab_9_8_port, B => CARRYB_8_8_port, CI => 
                           SUMB_8_9_port, CO => CARRYB_9_8_port, S => 
                           SUMB_9_8_port);
   S2_9_9 : FA_X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, CI => 
                           SUMB_8_10_port, CO => CARRYB_9_9_port, S => 
                           SUMB_9_9_port);
   S2_9_10 : FA_X1 port map( A => CARRYB_8_10_port, B => ab_9_10_port, CI => 
                           SUMB_8_11_port, CO => CARRYB_9_10_port, S => 
                           SUMB_9_10_port);
   S2_9_11 : FA_X1 port map( A => CARRYB_8_11_port, B => ab_9_11_port, CI => 
                           SUMB_8_12_port, CO => CARRYB_9_11_port, S => 
                           SUMB_9_11_port);
   S2_9_12 : FA_X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, CI => 
                           SUMB_8_13_port, CO => CARRYB_9_12_port, S => 
                           SUMB_9_12_port);
   S2_9_13 : FA_X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, CI => 
                           SUMB_8_14_port, CO => CARRYB_9_13_port, S => 
                           SUMB_9_13_port);
   S3_9_14 : FA_X1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, CI => 
                           ab_8_15_port, CO => CARRYB_9_14_port, S => 
                           SUMB_9_14_port);
   S1_8_0 : FA_X1 port map( A => ab_8_0_port, B => CARRYB_7_0_port, CI => 
                           SUMB_7_1_port, CO => CARRYB_8_0_port, S => A1_6_port
                           );
   S2_8_1 : FA_X1 port map( A => ab_8_1_port, B => CARRYB_7_1_port, CI => 
                           SUMB_7_2_port, CO => CARRYB_8_1_port, S => 
                           SUMB_8_1_port);
   S2_8_2 : FA_X1 port map( A => ab_8_2_port, B => CARRYB_7_2_port, CI => 
                           SUMB_7_3_port, CO => CARRYB_8_2_port, S => 
                           SUMB_8_2_port);
   S2_8_3 : FA_X1 port map( A => CARRYB_7_3_port, B => ab_8_3_port, CI => 
                           SUMB_7_4_port, CO => CARRYB_8_3_port, S => 
                           SUMB_8_3_port);
   S2_8_4 : FA_X1 port map( A => ab_8_4_port, B => CARRYB_7_4_port, CI => 
                           SUMB_7_5_port, CO => CARRYB_8_4_port, S => 
                           SUMB_8_4_port);
   S2_8_5 : FA_X1 port map( A => CARRYB_7_5_port, B => ab_8_5_port, CI => 
                           SUMB_7_6_port, CO => CARRYB_8_5_port, S => 
                           SUMB_8_5_port);
   S2_8_10 : FA_X1 port map( A => CARRYB_7_10_port, B => ab_8_10_port, CI => 
                           SUMB_7_11_port, CO => CARRYB_8_10_port, S => 
                           SUMB_8_10_port);
   S2_8_11 : FA_X1 port map( A => CARRYB_7_11_port, B => ab_8_11_port, CI => 
                           SUMB_7_12_port, CO => CARRYB_8_11_port, S => 
                           SUMB_8_11_port);
   S2_8_12 : FA_X1 port map( A => CARRYB_7_12_port, B => ab_8_12_port, CI => 
                           SUMB_7_13_port, CO => CARRYB_8_12_port, S => 
                           SUMB_8_12_port);
   S2_8_13 : FA_X1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, CI => 
                           SUMB_7_14_port, CO => CARRYB_8_13_port, S => 
                           SUMB_8_13_port);
   S3_8_14 : FA_X1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, CI => 
                           ab_7_15_port, CO => CARRYB_8_14_port, S => 
                           SUMB_8_14_port);
   S1_7_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => A1_5_port
                           );
   S2_7_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S2_7_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S2_7_3 : FA_X1 port map( A => CARRYB_6_3_port, B => ab_7_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S2_7_4 : FA_X1 port map( A => CARRYB_6_4_port, B => ab_7_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S2_7_5 : FA_X1 port map( A => CARRYB_6_5_port, B => ab_7_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S2_7_6 : FA_X1 port map( A => CARRYB_6_6_port, B => ab_7_6_port, CI => 
                           SUMB_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S2_7_10 : FA_X1 port map( A => ab_7_10_port, B => CARRYB_6_10_port, CI => 
                           SUMB_6_11_port, CO => CARRYB_7_10_port, S => 
                           SUMB_7_10_port);
   S2_7_11 : FA_X1 port map( A => CARRYB_6_11_port, B => ab_7_11_port, CI => 
                           SUMB_6_12_port, CO => CARRYB_7_11_port, S => 
                           SUMB_7_11_port);
   S2_7_12 : FA_X1 port map( A => CARRYB_6_12_port, B => ab_7_12_port, CI => 
                           SUMB_6_13_port, CO => CARRYB_7_12_port, S => 
                           SUMB_7_12_port);
   S2_7_13 : FA_X1 port map( A => SUMB_6_14_port, B => ab_7_13_port, CI => 
                           CARRYB_6_13_port, CO => CARRYB_7_13_port, S => 
                           SUMB_7_13_port);
   S3_7_14 : FA_X1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, CI => 
                           ab_6_15_port, CO => CARRYB_7_14_port, S => 
                           SUMB_7_14_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => CARRYB_5_5_port, B => ab_6_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S2_6_6 : FA_X1 port map( A => CARRYB_5_6_port, B => ab_6_6_port, CI => 
                           SUMB_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S2_6_7 : FA_X1 port map( A => CARRYB_5_7_port, B => ab_6_7_port, CI => 
                           SUMB_5_8_port, CO => CARRYB_6_7_port, S => 
                           SUMB_6_7_port);
   S2_6_11 : FA_X1 port map( A => ab_6_11_port, B => CARRYB_5_11_port, CI => 
                           SUMB_5_12_port, CO => CARRYB_6_11_port, S => 
                           SUMB_6_11_port);
   S2_6_12 : FA_X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, CI => 
                           SUMB_5_13_port, CO => CARRYB_6_12_port, S => 
                           SUMB_6_12_port);
   S2_6_13 : FA_X1 port map( A => CARRYB_5_13_port, B => ab_6_13_port, CI => 
                           SUMB_5_14_port, CO => CARRYB_6_13_port, S => 
                           SUMB_6_13_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => CARRYB_4_5_port, B => ab_5_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S2_5_6 : FA_X1 port map( A => CARRYB_4_6_port, B => ab_5_6_port, CI => 
                           SUMB_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S2_5_7 : FA_X1 port map( A => CARRYB_4_7_port, B => ab_5_7_port, CI => 
                           SUMB_4_8_port, CO => CARRYB_5_7_port, S => 
                           SUMB_5_7_port);
   S2_5_8 : FA_X1 port map( A => CARRYB_4_8_port, B => ab_5_8_port, CI => 
                           SUMB_4_9_port, CO => CARRYB_5_8_port, S => 
                           SUMB_5_8_port);
   S2_5_11 : FA_X1 port map( A => ab_5_11_port, B => CARRYB_4_11_port, CI => 
                           SUMB_4_12_port, CO => CARRYB_5_11_port, S => 
                           SUMB_5_11_port);
   S2_5_12 : FA_X1 port map( A => CARRYB_4_12_port, B => ab_5_12_port, CI => 
                           SUMB_4_13_port, CO => CARRYB_5_12_port, S => 
                           SUMB_5_12_port);
   S2_5_13 : FA_X1 port map( A => CARRYB_4_13_port, B => ab_5_13_port, CI => 
                           SUMB_4_14_port, CO => CARRYB_5_13_port, S => 
                           SUMB_5_13_port);
   S3_5_14 : FA_X1 port map( A => ab_5_14_port, B => CARRYB_4_14_port, CI => 
                           ab_4_15_port, CO => CARRYB_5_14_port, S => 
                           SUMB_5_14_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => CARRYB_3_3_port, B => ab_4_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S2_4_6 : FA_X1 port map( A => CARRYB_3_6_port, B => ab_4_6_port, CI => 
                           SUMB_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S2_4_7 : FA_X1 port map( A => CARRYB_3_7_port, B => ab_4_7_port, CI => 
                           SUMB_3_8_port, CO => CARRYB_4_7_port, S => 
                           SUMB_4_7_port);
   S2_4_8 : FA_X1 port map( A => ab_4_8_port, B => CARRYB_3_8_port, CI => 
                           SUMB_3_9_port, CO => CARRYB_4_8_port, S => 
                           SUMB_4_8_port);
   S2_4_9 : FA_X1 port map( A => CARRYB_3_9_port, B => ab_4_9_port, CI => 
                           SUMB_3_10_port, CO => CARRYB_4_9_port, S => 
                           SUMB_4_9_port);
   S2_4_13 : FA_X1 port map( A => ab_4_13_port, B => SUMB_3_14_port, CI => 
                           CARRYB_3_13_port, CO => CARRYB_4_13_port, S => 
                           SUMB_4_13_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S2_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           SUMB_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S2_3_7 : FA_X1 port map( A => CARRYB_2_7_port, B => ab_3_7_port, CI => 
                           SUMB_2_8_port, CO => CARRYB_3_7_port, S => 
                           SUMB_3_7_port);
   S2_3_8 : FA_X1 port map( A => ab_3_8_port, B => CARRYB_2_8_port, CI => 
                           SUMB_2_9_port, CO => CARRYB_3_8_port, S => 
                           SUMB_3_8_port);
   S2_3_9 : FA_X1 port map( A => ab_3_9_port, B => CARRYB_2_9_port, CI => 
                           SUMB_2_10_port, CO => CARRYB_3_9_port, S => 
                           SUMB_3_9_port);
   S2_3_10 : FA_X1 port map( A => CARRYB_2_10_port, B => ab_3_10_port, CI => 
                           SUMB_2_11_port, CO => CARRYB_3_10_port, S => 
                           SUMB_3_10_port);
   S2_3_13 : FA_X1 port map( A => ab_3_13_port, B => CARRYB_2_13_port, CI => 
                           SUMB_2_14_port, CO => CARRYB_3_13_port, S => 
                           SUMB_3_13_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n4, CI => n20, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n19, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n18, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n3, CI => n30, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n16, CI => n29, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n15, CI => n28, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S2_2_7 : FA_X1 port map( A => ab_2_7_port, B => n13, CI => n22, CO => 
                           CARRYB_2_7_port, S => SUMB_2_7_port);
   S2_2_8 : FA_X1 port map( A => ab_2_8_port, B => n8, CI => n24, CO => 
                           CARRYB_2_8_port, S => SUMB_2_8_port);
   S2_2_10 : FA_X1 port map( A => n7, B => ab_2_10_port, CI => n23, CO => 
                           CARRYB_2_10_port, S => SUMB_2_10_port);
   S2_2_11 : FA_X1 port map( A => ab_2_11_port, B => n9, CI => n25, CO => 
                           CARRYB_2_11_port, S => SUMB_2_11_port);
   U18 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n19);
   U19 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n20);
   U26 : XOR2_X1 port map( A => ab_1_7_port, B => ab_0_8_port, Z => n27);
   U28 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n29);
   U29 : XOR2_X1 port map( A => n292, B => ab_0_5_port, Z => n30);
   U32 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U37 : XOR2_X1 port map( A => CARRYB_15_5_port, B => SUMB_15_6_port, Z => n36
                           );
   U38 : XOR2_X1 port map( A => CARRYB_15_7_port, B => SUMB_15_8_port, Z => n37
                           );
   U39 : XOR2_X1 port map( A => CARRYB_15_9_port, B => SUMB_15_10_port, Z => 
                           n38);
   U40 : XOR2_X1 port map( A => CARRYB_15_11_port, B => SUMB_15_12_port, Z => 
                           n39);
   U41 : XOR2_X1 port map( A => CARRYB_15_13_port, B => SUMB_15_14_port, Z => 
                           n40);
   U52 : XOR2_X1 port map( A => CARRYB_15_6_port, B => SUMB_15_7_port, Z => n51
                           );
   U53 : XOR2_X1 port map( A => CARRYB_15_8_port, B => SUMB_15_9_port, Z => n52
                           );
   U54 : XOR2_X1 port map( A => CARRYB_15_10_port, B => SUMB_15_11_port, Z => 
                           n53);
   U55 : XOR2_X1 port map( A => CARRYB_15_12_port, B => SUMB_15_13_port, Z => 
                           n54);
   U63 : XOR2_X1 port map( A => CARRYB_15_14_port, B => SUMB_15_15_port, Z => 
                           n62);
   U97 : XOR2_X1 port map( A => CARRYB_15_15_port, B => n125, Z => n63);
   U98 : NOR2_X1 port map( A1 => net74673, A2 => n184, ZN => ab_9_9_port);
   U99 : NOR2_X1 port map( A1 => net74673, A2 => n192, ZN => ab_9_8_port);
   U101 : NOR2_X1 port map( A1 => net74673, A2 => n189, ZN => ab_9_6_port);
   U102 : NOR2_X1 port map( A1 => net74673, A2 => n186, ZN => ab_9_5_port);
   U103 : NOR2_X1 port map( A1 => net74673, A2 => n248, ZN => ab_9_4_port);
   U104 : NOR2_X1 port map( A1 => net74673, A2 => n278, ZN => ab_9_3_port);
   U105 : NOR2_X1 port map( A1 => net74673, A2 => n181, ZN => ab_9_2_port);
   U106 : NOR2_X1 port map( A1 => net74673, A2 => n280, ZN => ab_9_1_port);
   U108 : NOR2_X1 port map( A1 => net74673, A2 => net82535, ZN => ab_9_14_port)
                           ;
   U109 : NOR2_X1 port map( A1 => net74673, A2 => net118627, ZN => ab_9_13_port
                           );
   U110 : NOR2_X1 port map( A1 => net74673, A2 => net97008, ZN => ab_9_12_port)
                           ;
   U111 : NOR2_X1 port map( A1 => net74673, A2 => net82653, ZN => ab_9_11_port)
                           ;
   U112 : NOR2_X1 port map( A1 => net74673, A2 => net82724, ZN => ab_9_10_port)
                           ;
   U113 : NOR2_X1 port map( A1 => net74673, A2 => net74680, ZN => ab_9_0_port);
   U114 : NOR2_X1 port map( A1 => n184, A2 => n287, ZN => ab_8_9_port);
   U115 : NOR2_X1 port map( A1 => n192, A2 => n287, ZN => ab_8_8_port);
   U116 : NOR2_X1 port map( A1 => net82987, A2 => n287, ZN => ab_8_7_port);
   U117 : NOR2_X1 port map( A1 => n189, A2 => n287, ZN => ab_8_6_port);
   U118 : NOR2_X1 port map( A1 => n186, A2 => n287, ZN => ab_8_5_port);
   U119 : NOR2_X1 port map( A1 => n248, A2 => n287, ZN => ab_8_4_port);
   U120 : NOR2_X1 port map( A1 => n278, A2 => n287, ZN => ab_8_3_port);
   U121 : NOR2_X1 port map( A1 => n181, A2 => n287, ZN => ab_8_2_port);
   U122 : NOR2_X1 port map( A1 => n280, A2 => n287, ZN => ab_8_1_port);
   U124 : NOR2_X1 port map( A1 => net82535, A2 => n287, ZN => ab_8_14_port);
   U125 : NOR2_X1 port map( A1 => net118627, A2 => n287, ZN => ab_8_13_port);
   U126 : NOR2_X1 port map( A1 => net97008, A2 => n287, ZN => ab_8_12_port);
   U127 : NOR2_X1 port map( A1 => net82653, A2 => n287, ZN => ab_8_11_port);
   U128 : NOR2_X1 port map( A1 => net82724, A2 => n287, ZN => ab_8_10_port);
   U129 : NOR2_X1 port map( A1 => net74680, A2 => n287, ZN => ab_8_0_port);
   U130 : NOR2_X1 port map( A1 => n184, A2 => n288, ZN => ab_7_9_port);
   U131 : NOR2_X1 port map( A1 => n192, A2 => n288, ZN => ab_7_8_port);
   U132 : NOR2_X1 port map( A1 => net82987, A2 => n288, ZN => ab_7_7_port);
   U133 : NOR2_X1 port map( A1 => n189, A2 => n288, ZN => ab_7_6_port);
   U134 : NOR2_X1 port map( A1 => n186, A2 => n288, ZN => ab_7_5_port);
   U135 : NOR2_X1 port map( A1 => n248, A2 => n288, ZN => ab_7_4_port);
   U136 : NOR2_X1 port map( A1 => n278, A2 => n288, ZN => ab_7_3_port);
   U137 : NOR2_X1 port map( A1 => n181, A2 => n288, ZN => ab_7_2_port);
   U138 : NOR2_X1 port map( A1 => n280, A2 => n288, ZN => ab_7_1_port);
   U140 : NOR2_X1 port map( A1 => net82535, A2 => n288, ZN => ab_7_14_port);
   U141 : NOR2_X1 port map( A1 => net118627, A2 => n288, ZN => ab_7_13_port);
   U142 : NOR2_X1 port map( A1 => net97008, A2 => n288, ZN => ab_7_12_port);
   U143 : NOR2_X1 port map( A1 => net82653, A2 => n288, ZN => ab_7_11_port);
   U144 : NOR2_X1 port map( A1 => net82724, A2 => n288, ZN => ab_7_10_port);
   U145 : NOR2_X1 port map( A1 => net74680, A2 => n288, ZN => ab_7_0_port);
   U146 : NOR2_X1 port map( A1 => n184, A2 => n265, ZN => ab_6_9_port);
   U147 : NOR2_X1 port map( A1 => n192, A2 => n266, ZN => ab_6_8_port);
   U148 : NOR2_X1 port map( A1 => net82987, A2 => n265, ZN => ab_6_7_port);
   U149 : NOR2_X1 port map( A1 => n189, A2 => n266, ZN => ab_6_6_port);
   U150 : NOR2_X1 port map( A1 => n186, A2 => n265, ZN => ab_6_5_port);
   U151 : NOR2_X1 port map( A1 => n248, A2 => n266, ZN => ab_6_4_port);
   U152 : NOR2_X1 port map( A1 => n278, A2 => n265, ZN => ab_6_3_port);
   U153 : NOR2_X1 port map( A1 => n181, A2 => n266, ZN => ab_6_2_port);
   U154 : NOR2_X1 port map( A1 => n280, A2 => n265, ZN => ab_6_1_port);
   U156 : NOR2_X1 port map( A1 => net82535, A2 => n266, ZN => ab_6_14_port);
   U157 : NOR2_X1 port map( A1 => net118627, A2 => n265, ZN => ab_6_13_port);
   U158 : NOR2_X1 port map( A1 => net97008, A2 => n266, ZN => ab_6_12_port);
   U159 : NOR2_X1 port map( A1 => net82653, A2 => n289, ZN => ab_6_11_port);
   U160 : NOR2_X1 port map( A1 => net82724, A2 => n265, ZN => ab_6_10_port);
   U161 : NOR2_X1 port map( A1 => net74680, A2 => n289, ZN => ab_6_0_port);
   U162 : NOR2_X1 port map( A1 => n184, A2 => net74669, ZN => ab_5_9_port);
   U163 : NOR2_X1 port map( A1 => n192, A2 => net74669, ZN => ab_5_8_port);
   U164 : NOR2_X1 port map( A1 => net82987, A2 => net74669, ZN => ab_5_7_port);
   U165 : NOR2_X1 port map( A1 => n189, A2 => net74669, ZN => ab_5_6_port);
   U166 : NOR2_X1 port map( A1 => n186, A2 => net74669, ZN => ab_5_5_port);
   U167 : NOR2_X1 port map( A1 => n248, A2 => net74669, ZN => ab_5_4_port);
   U168 : NOR2_X1 port map( A1 => n278, A2 => net74669, ZN => ab_5_3_port);
   U169 : NOR2_X1 port map( A1 => n181, A2 => net74669, ZN => ab_5_2_port);
   U170 : NOR2_X1 port map( A1 => n280, A2 => net74669, ZN => ab_5_1_port);
   U172 : NOR2_X1 port map( A1 => net82535, A2 => net74669, ZN => ab_5_14_port)
                           ;
   U173 : NOR2_X1 port map( A1 => net118627, A2 => net74669, ZN => ab_5_13_port
                           );
   U174 : NOR2_X1 port map( A1 => net97008, A2 => net74669, ZN => ab_5_12_port)
                           ;
   U178 : NOR2_X1 port map( A1 => n184, A2 => n290, ZN => ab_4_9_port);
   U179 : NOR2_X1 port map( A1 => n274, A2 => n290, ZN => ab_4_8_port);
   U180 : NOR2_X1 port map( A1 => net82987, A2 => n290, ZN => ab_4_7_port);
   U181 : NOR2_X1 port map( A1 => n189, A2 => n290, ZN => ab_4_6_port);
   U182 : NOR2_X1 port map( A1 => n186, A2 => n290, ZN => ab_4_5_port);
   U183 : NOR2_X1 port map( A1 => n248, A2 => n290, ZN => ab_4_4_port);
   U184 : NOR2_X1 port map( A1 => n278, A2 => n290, ZN => ab_4_3_port);
   U185 : NOR2_X1 port map( A1 => n181, A2 => n290, ZN => ab_4_2_port);
   U186 : NOR2_X1 port map( A1 => n280, A2 => n290, ZN => ab_4_1_port);
   U188 : NOR2_X1 port map( A1 => net74694, A2 => n290, ZN => ab_4_14_port);
   U189 : NOR2_X1 port map( A1 => net118627, A2 => n290, ZN => ab_4_13_port);
   U190 : NOR2_X1 port map( A1 => n290, A2 => net97008, ZN => ab_4_12_port);
   U191 : NOR2_X1 port map( A1 => net82653, A2 => n290, ZN => ab_4_11_port);
   U192 : NOR2_X1 port map( A1 => net82724, A2 => n290, ZN => ab_4_10_port);
   U193 : NOR2_X1 port map( A1 => net74680, A2 => n290, ZN => ab_4_0_port);
   U194 : NOR2_X1 port map( A1 => n184, A2 => net82975, ZN => ab_3_9_port);
   U195 : NOR2_X1 port map( A1 => n274, A2 => net82976, ZN => ab_3_8_port);
   U196 : NOR2_X1 port map( A1 => net82987, A2 => net82976, ZN => ab_3_7_port);
   U197 : NOR2_X1 port map( A1 => n189, A2 => net82975, ZN => ab_3_6_port);
   U198 : NOR2_X1 port map( A1 => n186, A2 => net82976, ZN => ab_3_5_port);
   U199 : NOR2_X1 port map( A1 => n248, A2 => net82976, ZN => ab_3_4_port);
   U200 : NOR2_X1 port map( A1 => n278, A2 => net82976, ZN => ab_3_3_port);
   U201 : NOR2_X1 port map( A1 => n181, A2 => net82975, ZN => ab_3_2_port);
   U202 : NOR2_X1 port map( A1 => n280, A2 => net82976, ZN => ab_3_1_port);
   U205 : NOR2_X1 port map( A1 => net118627, A2 => net82975, ZN => ab_3_13_port
                           );
   U208 : NOR2_X1 port map( A1 => net82724, A2 => net82976, ZN => ab_3_10_port)
                           ;
   U209 : NOR2_X1 port map( A1 => net74680, A2 => net82975, ZN => ab_3_0_port);
   U210 : NOR2_X1 port map( A1 => n243, A2 => net83102, ZN => ab_2_9_port);
   U211 : NOR2_X1 port map( A1 => n274, A2 => net83102, ZN => ab_2_8_port);
   U213 : NOR2_X1 port map( A1 => n275, A2 => net74666, ZN => ab_2_6_port);
   U214 : NOR2_X1 port map( A1 => n276, A2 => net74666, ZN => ab_2_5_port);
   U215 : NOR2_X1 port map( A1 => n187, A2 => net83102, ZN => ab_2_4_port);
   U216 : NOR2_X1 port map( A1 => n278, A2 => net83102, ZN => ab_2_3_port);
   U217 : NOR2_X1 port map( A1 => n181, A2 => net83102, ZN => ab_2_2_port);
   U218 : NOR2_X1 port map( A1 => n280, A2 => net83102, ZN => ab_2_1_port);
   U220 : NOR2_X1 port map( A1 => net74694, A2 => net83102, ZN => ab_2_14_port)
                           ;
   U221 : NOR2_X1 port map( A1 => net74693, A2 => net83102, ZN => ab_2_13_port)
                           ;
   U223 : NOR2_X1 port map( A1 => net74666, A2 => net74691, ZN => ab_2_11_port)
                           ;
   U224 : NOR2_X1 port map( A1 => net74666, A2 => net74690, ZN => ab_2_10_port)
                           ;
   U225 : NOR2_X1 port map( A1 => net74680, A2 => net83102, ZN => ab_2_0_port);
   U229 : NOR2_X1 port map( A1 => n275, A2 => net77076, ZN => ab_1_6_port);
   U230 : NOR2_X1 port map( A1 => n276, A2 => net77076, ZN => ab_1_5_port);
   U234 : NOR2_X1 port map( A1 => n280, A2 => net77076, ZN => ab_1_1_port);
   U241 : NOR2_X1 port map( A1 => net74680, A2 => net77076, ZN => ab_1_0_port);
   U251 : NOR2_X1 port map( A1 => n272, A2 => n281, ZN => ab_15_15_port);
   U258 : NOR2_X1 port map( A1 => n281, A2 => n125, ZN => n99);
   U259 : NOR2_X1 port map( A1 => n184, A2 => n282, ZN => ab_14_9_port);
   U260 : NOR2_X1 port map( A1 => n192, A2 => n282, ZN => ab_14_8_port);
   U261 : NOR2_X1 port map( A1 => net82987, A2 => n282, ZN => ab_14_7_port);
   U262 : NOR2_X1 port map( A1 => n189, A2 => n282, ZN => ab_14_6_port);
   U263 : NOR2_X1 port map( A1 => n186, A2 => n282, ZN => ab_14_5_port);
   U264 : NOR2_X1 port map( A1 => n248, A2 => n282, ZN => ab_14_4_port);
   U265 : NOR2_X1 port map( A1 => n278, A2 => n282, ZN => ab_14_3_port);
   U266 : NOR2_X1 port map( A1 => n181, A2 => n282, ZN => ab_14_2_port);
   U267 : NOR2_X1 port map( A1 => n280, A2 => n282, ZN => ab_14_1_port);
   U269 : NOR2_X1 port map( A1 => net82535, A2 => n282, ZN => ab_14_14_port);
   U270 : NOR2_X1 port map( A1 => net118627, A2 => n282, ZN => ab_14_13_port);
   U271 : NOR2_X1 port map( A1 => net97008, A2 => n282, ZN => ab_14_12_port);
   U272 : NOR2_X1 port map( A1 => net82653, A2 => n282, ZN => ab_14_11_port);
   U273 : NOR2_X1 port map( A1 => net82724, A2 => n282, ZN => ab_14_10_port);
   U274 : NOR2_X1 port map( A1 => net74680, A2 => n282, ZN => ab_14_0_port);
   U275 : NOR2_X1 port map( A1 => n184, A2 => n283, ZN => ab_13_9_port);
   U276 : NOR2_X1 port map( A1 => n192, A2 => n283, ZN => ab_13_8_port);
   U277 : NOR2_X1 port map( A1 => net82987, A2 => n283, ZN => ab_13_7_port);
   U278 : NOR2_X1 port map( A1 => n189, A2 => n283, ZN => ab_13_6_port);
   U279 : NOR2_X1 port map( A1 => n186, A2 => n283, ZN => ab_13_5_port);
   U280 : NOR2_X1 port map( A1 => n248, A2 => n283, ZN => ab_13_4_port);
   U281 : NOR2_X1 port map( A1 => n278, A2 => n283, ZN => ab_13_3_port);
   U282 : NOR2_X1 port map( A1 => n181, A2 => n283, ZN => ab_13_2_port);
   U283 : NOR2_X1 port map( A1 => n280, A2 => n283, ZN => ab_13_1_port);
   U285 : NOR2_X1 port map( A1 => net82535, A2 => n283, ZN => ab_13_14_port);
   U286 : NOR2_X1 port map( A1 => net118627, A2 => n283, ZN => ab_13_13_port);
   U287 : NOR2_X1 port map( A1 => net97008, A2 => n283, ZN => ab_13_12_port);
   U288 : NOR2_X1 port map( A1 => net82653, A2 => n283, ZN => ab_13_11_port);
   U289 : NOR2_X1 port map( A1 => net82724, A2 => n283, ZN => ab_13_10_port);
   U290 : NOR2_X1 port map( A1 => net74680, A2 => n283, ZN => ab_13_0_port);
   U291 : NOR2_X1 port map( A1 => n184, A2 => n284, ZN => ab_12_9_port);
   U292 : NOR2_X1 port map( A1 => n192, A2 => n284, ZN => ab_12_8_port);
   U293 : NOR2_X1 port map( A1 => net82987, A2 => n284, ZN => ab_12_7_port);
   U294 : NOR2_X1 port map( A1 => n189, A2 => n284, ZN => ab_12_6_port);
   U295 : NOR2_X1 port map( A1 => n186, A2 => n284, ZN => ab_12_5_port);
   U296 : NOR2_X1 port map( A1 => n248, A2 => n284, ZN => ab_12_4_port);
   U297 : NOR2_X1 port map( A1 => n278, A2 => n284, ZN => ab_12_3_port);
   U298 : NOR2_X1 port map( A1 => n181, A2 => n284, ZN => ab_12_2_port);
   U299 : NOR2_X1 port map( A1 => n280, A2 => n284, ZN => ab_12_1_port);
   U301 : NOR2_X1 port map( A1 => net82535, A2 => n284, ZN => ab_12_14_port);
   U302 : NOR2_X1 port map( A1 => net118627, A2 => n284, ZN => ab_12_13_port);
   U303 : NOR2_X1 port map( A1 => net97008, A2 => n284, ZN => ab_12_12_port);
   U304 : NOR2_X1 port map( A1 => net82653, A2 => n284, ZN => ab_12_11_port);
   U305 : NOR2_X1 port map( A1 => net82724, A2 => n284, ZN => ab_12_10_port);
   U306 : NOR2_X1 port map( A1 => net74680, A2 => n284, ZN => ab_12_0_port);
   U307 : NOR2_X1 port map( A1 => n184, A2 => n285, ZN => ab_11_9_port);
   U308 : NOR2_X1 port map( A1 => n192, A2 => n285, ZN => ab_11_8_port);
   U309 : NOR2_X1 port map( A1 => net82987, A2 => n285, ZN => ab_11_7_port);
   U310 : NOR2_X1 port map( A1 => n189, A2 => n285, ZN => ab_11_6_port);
   U311 : NOR2_X1 port map( A1 => n186, A2 => n285, ZN => ab_11_5_port);
   U312 : NOR2_X1 port map( A1 => n248, A2 => n285, ZN => ab_11_4_port);
   U313 : NOR2_X1 port map( A1 => n278, A2 => n285, ZN => ab_11_3_port);
   U314 : NOR2_X1 port map( A1 => n181, A2 => n285, ZN => ab_11_2_port);
   U315 : NOR2_X1 port map( A1 => n280, A2 => n285, ZN => ab_11_1_port);
   U317 : NOR2_X1 port map( A1 => net82535, A2 => n285, ZN => ab_11_14_port);
   U318 : NOR2_X1 port map( A1 => net118627, A2 => n285, ZN => ab_11_13_port);
   U319 : NOR2_X1 port map( A1 => net97008, A2 => n285, ZN => ab_11_12_port);
   U320 : NOR2_X1 port map( A1 => net82653, A2 => n285, ZN => ab_11_11_port);
   U321 : NOR2_X1 port map( A1 => net82724, A2 => n285, ZN => ab_11_10_port);
   U322 : NOR2_X1 port map( A1 => net74680, A2 => n285, ZN => ab_11_0_port);
   U323 : NOR2_X1 port map( A1 => n184, A2 => n286, ZN => ab_10_9_port);
   U324 : NOR2_X1 port map( A1 => n192, A2 => n286, ZN => ab_10_8_port);
   U325 : NOR2_X1 port map( A1 => net82987, A2 => n286, ZN => ab_10_7_port);
   U326 : NOR2_X1 port map( A1 => n189, A2 => n286, ZN => ab_10_6_port);
   U327 : NOR2_X1 port map( A1 => n186, A2 => n286, ZN => ab_10_5_port);
   U328 : NOR2_X1 port map( A1 => n248, A2 => n286, ZN => ab_10_4_port);
   U329 : NOR2_X1 port map( A1 => n278, A2 => n286, ZN => ab_10_3_port);
   U330 : NOR2_X1 port map( A1 => n181, A2 => n286, ZN => ab_10_2_port);
   U331 : NOR2_X1 port map( A1 => n280, A2 => n286, ZN => ab_10_1_port);
   U333 : NOR2_X1 port map( A1 => net82535, A2 => n286, ZN => ab_10_14_port);
   U334 : NOR2_X1 port map( A1 => net118627, A2 => n286, ZN => ab_10_13_port);
   U335 : NOR2_X1 port map( A1 => net97008, A2 => n286, ZN => ab_10_12_port);
   U336 : NOR2_X1 port map( A1 => net82653, A2 => n286, ZN => ab_10_11_port);
   U337 : NOR2_X1 port map( A1 => net82724, A2 => n286, ZN => ab_10_10_port);
   U338 : NOR2_X1 port map( A1 => net74680, A2 => n286, ZN => ab_10_0_port);
   U339 : NOR2_X1 port map( A1 => n243, A2 => net77069, ZN => ab_0_9_port);
   U340 : NOR2_X1 port map( A1 => n274, A2 => net77069, ZN => ab_0_8_port);
   U342 : NOR2_X1 port map( A1 => n275, A2 => net77069, ZN => ab_0_6_port);
   U343 : NOR2_X1 port map( A1 => n276, A2 => net83062, ZN => ab_0_5_port);
   U344 : NOR2_X1 port map( A1 => n187, A2 => net83062, ZN => ab_0_4_port);
   U345 : NOR2_X1 port map( A1 => n278, A2 => net83062, ZN => ab_0_3_port);
   U346 : NOR2_X1 port map( A1 => n181, A2 => net83062, ZN => ab_0_2_port);
   U347 : NOR2_X1 port map( A1 => n280, A2 => net77069, ZN => ab_0_1_port);
   U349 : NOR2_X1 port map( A1 => n141, A2 => TC, ZN => n98);
   U354 : NOR2_X1 port map( A1 => net74690, A2 => net77069, ZN => ab_0_10_port)
                           ;
   U355 : NOR2_X1 port map( A1 => B(15), A2 => n291, ZN => QB);
   U356 : NOR2_X1 port map( A1 => A(15), A2 => n291, ZN => QA);
   U357 : NOR2_X1 port map( A1 => net74680, A2 => net77069, ZN => PRODUCT(0));
   U34 : NOR2_X1 port map( A1 => n281, A2 => n291, ZN => ZA);
   n100 <= '0';
   n101 <= '0';
   U177 : NOR2_X1 port map( A1 => net74680, A2 => net74669, ZN => ab_5_0_port);
   U175 : NOR2_X1 port map( A1 => net82653, A2 => net74669, ZN => ab_5_11_port)
                           ;
   U176 : NOR2_X1 port map( A1 => net82724, A2 => net74669, ZN => ab_5_10_port)
                           ;
   S2_13_2 : FA_X1 port map( A => CARRYB_12_2_port, B => ab_13_2_port, CI => 
                           SUMB_12_3_port, CO => CARRYB_13_2_port, S => 
                           SUMB_13_2_port);
   S2_12_2 : FA_X1 port map( A => CARRYB_11_2_port, B => ab_12_2_port, CI => 
                           SUMB_11_3_port, CO => CARRYB_12_2_port, S => 
                           SUMB_12_2_port);
   S2_12_3 : FA_X1 port map( A => CARRYB_11_3_port, B => ab_12_3_port, CI => 
                           SUMB_11_4_port, CO => CARRYB_12_3_port, S => 
                           SUMB_12_3_port);
   S4_1 : FA_X1 port map( A => CARRYB_14_1_port, B => ab_15_1_port, CI => 
                           SUMB_14_2_port, CO => CARRYB_15_1_port, S => 
                           SUMB_15_1_port);
   S4_2 : FA_X1 port map( A => ab_15_2_port, B => CARRYB_14_2_port, CI => 
                           SUMB_14_3_port, CO => CARRYB_15_2_port, S => 
                           SUMB_15_2_port);
   U212 : NOR2_X1 port map( A1 => net74687, A2 => net83102, ZN => ab_2_7_port);
   U341 : NOR2_X1 port map( A1 => net74687, A2 => net77069, ZN => ab_0_7_port);
   U100 : NOR2_X1 port map( A1 => net74673, A2 => net82987, ZN => ab_9_7_port);
   S2_9_7 : FA_X1 port map( A => CARRYB_8_7_port, B => ab_9_7_port, CI => 
                           SUMB_8_8_port, CO => CARRYB_9_7_port, S => 
                           SUMB_9_7_port);
   S2_10_6 : FA_X1 port map( A => ab_10_6_port, B => CARRYB_9_6_port, CI => 
                           SUMB_9_7_port, CO => CARRYB_10_6_port, S => 
                           SUMB_10_6_port);
   S2_11_5 : FA_X1 port map( A => CARRYB_10_5_port, B => ab_11_5_port, CI => 
                           SUMB_10_6_port, CO => CARRYB_11_5_port, S => 
                           SUMB_11_5_port);
   S2_12_4 : FA_X1 port map( A => ab_12_4_port, B => CARRYB_11_4_port, CI => 
                           SUMB_11_5_port, CO => CARRYB_12_4_port, S => 
                           SUMB_12_4_port);
   S2_14_2 : FA_X1 port map( A => ab_14_2_port, B => CARRYB_13_2_port, CI => 
                           SUMB_13_3_port, CO => CARRYB_14_2_port, S => 
                           SUMB_14_2_port);
   S2_13_3 : FA_X1 port map( A => CARRYB_12_3_port, B => ab_13_3_port, CI => 
                           SUMB_12_4_port, CO => CARRYB_13_3_port, S => 
                           SUMB_13_3_port);
   S2_11_3 : FA_X1 port map( A => CARRYB_10_3_port, B => ab_11_3_port, CI => 
                           SUMB_10_4_port, CO => CARRYB_11_3_port, S => 
                           SUMB_11_3_port);
   S2_11_4 : FA_X1 port map( A => CARRYB_10_4_port, B => ab_11_4_port, CI => 
                           SUMB_10_5_port, CO => CARRYB_11_4_port, S => 
                           SUMB_11_4_port);
   S2_10_4 : FA_X1 port map( A => CARRYB_9_4_port, B => ab_10_4_port, CI => 
                           SUMB_9_5_port, CO => CARRYB_10_4_port, S => 
                           SUMB_10_4_port);
   S2_10_5 : FA_X1 port map( A => CARRYB_9_5_port, B => ab_10_5_port, CI => 
                           SUMB_9_6_port, CO => CARRYB_10_5_port, S => 
                           SUMB_10_5_port);
   S2_9_5 : FA_X1 port map( A => CARRYB_8_5_port, B => ab_9_5_port, CI => 
                           SUMB_8_6_port, CO => CARRYB_9_5_port, S => 
                           SUMB_9_5_port);
   S2_9_6 : FA_X1 port map( A => CARRYB_8_6_port, B => ab_9_6_port, CI => 
                           SUMB_8_7_port, CO => CARRYB_9_6_port, S => 
                           SUMB_9_6_port);
   S2_8_6 : FA_X1 port map( A => CARRYB_7_6_port, B => ab_8_6_port, CI => 
                           SUMB_7_7_port, CO => CARRYB_8_6_port, S => 
                           SUMB_8_6_port);
   S2_8_7 : FA_X1 port map( A => CARRYB_7_7_port, B => ab_8_7_port, CI => 
                           SUMB_7_8_port, CO => CARRYB_8_7_port, S => 
                           SUMB_8_7_port);
   S2_7_7 : FA_X1 port map( A => CARRYB_6_7_port, B => ab_7_7_port, CI => 
                           SUMB_6_8_port, CO => CARRYB_7_7_port, S => 
                           SUMB_7_7_port);
   S2_7_8 : FA_X1 port map( A => CARRYB_6_8_port, B => ab_7_8_port, CI => 
                           SUMB_6_9_port, CO => CARRYB_7_8_port, S => 
                           SUMB_7_8_port);
   S2_6_8 : FA_X1 port map( A => CARRYB_5_8_port, B => ab_6_8_port, CI => 
                           SUMB_5_9_port, CO => CARRYB_6_8_port, S => 
                           SUMB_6_8_port);
   S2_6_9 : FA_X1 port map( A => CARRYB_5_9_port, B => ab_6_9_port, CI => 
                           SUMB_5_10_port, CO => CARRYB_6_9_port, S => 
                           SUMB_6_9_port);
   S2_5_9 : FA_X1 port map( A => CARRYB_4_9_port, B => ab_5_9_port, CI => 
                           SUMB_4_10_port, CO => CARRYB_5_9_port, S => 
                           SUMB_5_9_port);
   S2_5_10 : FA_X1 port map( A => CARRYB_4_10_port, B => ab_5_10_port, CI => 
                           SUMB_4_11_port, CO => CARRYB_5_10_port, S => 
                           SUMB_5_10_port);
   U353 : NOR2_X1 port map( A1 => net74691, A2 => net77069, ZN => ab_0_11_port)
                           ;
   U204 : NOR2_X1 port map( A1 => net74694, A2 => net82976, ZN => ab_3_14_port)
                           ;
   U207 : NOR2_X1 port map( A1 => net82653, A2 => net82975, ZN => ab_3_11_port)
                           ;
   U206 : NOR2_X1 port map( A1 => net82976, A2 => net74692, ZN => ab_3_12_port)
                           ;
   U222 : NOR2_X1 port map( A1 => net74666, A2 => net74692, ZN => ab_2_12_port)
                           ;
   S2_2_12 : FA_X1 port map( A => n11, B => ab_2_12_port, CI => n26, CO => 
                           CARRYB_2_12_port, S => SUMB_2_12_port);
   S2_4_10 : FA_X1 port map( A => CARRYB_3_10_port, B => ab_4_10_port, CI => 
                           SUMB_3_11_port, CO => CARRYB_4_10_port, S => 
                           SUMB_4_10_port);
   S2_3_11 : FA_X1 port map( A => CARRYB_2_11_port, B => ab_3_11_port, CI => 
                           SUMB_2_12_port, CO => CARRYB_3_11_port, S => 
                           SUMB_3_11_port);
   U23 : XNOR2_X1 port map( A => n105, B => SUMB_11_6_port, ZN => 
                           SUMB_12_5_port);
   U24 : XNOR2_X1 port map( A => ab_12_5_port, B => CARRYB_11_5_port, ZN => 
                           n105);
   U35 : XNOR2_X1 port map( A => net82534, B => net82716, ZN => n26);
   U50 : INV_X1 port map( A => B(14), ZN => net74694);
   U51 : INV_X1 port map( A => A(0), ZN => net74664);
   U67 : XNOR2_X1 port map( A => CARRYB_3_11_port, B => ab_4_11_port, ZN => 
                           net82396);
   U68 : XNOR2_X1 port map( A => ab_3_12_port, B => CARRYB_2_12_port, ZN => 
                           net82414);
   U69 : NAND2_X1 port map( A1 => SUMB_2_13_port, A2 => CARRYB_2_12_port, ZN =>
                           net82387);
   U70 : NAND2_X1 port map( A1 => ab_3_12_port, A2 => CARRYB_2_12_port, ZN => 
                           net82385);
   U71 : NAND2_X1 port map( A1 => A(1), A2 => B(13), ZN => net82716);
   U72 : NAND2_X1 port map( A1 => n102, A2 => B(12), ZN => net82986);
   U76 : INV_X1 port map( A => A(2), ZN => net74666);
   U78 : INV_X1 port map( A => B(12), ZN => net74692);
   U79 : CLKBUF_X1 port map( A => net74692, Z => net97008);
   U82 : INV_X1 port map( A => net74691, ZN => net82651);
   U83 : NAND2_X1 port map( A1 => net82651, A2 => net83064, ZN => net82980);
   U84 : INV_X1 port map( A => B(11), ZN => net74691);
   U85 : XNOR2_X1 port map( A => CARRYB_13_3_port, B => ab_14_3_port, ZN => 
                           net82608);
   U86 : NAND2_X1 port map( A1 => CARRYB_13_3_port, A2 => ab_14_3_port, ZN => 
                           net82597);
   U87 : NAND2_X1 port map( A1 => net82876, A2 => CARRYB_13_3_port, ZN => 
                           net82595);
   U88 : XNOR2_X1 port map( A => CARRYB_12_4_port, B => ab_13_4_port, ZN => 
                           net82778);
   U89 : NAND2_X1 port map( A1 => CARRYB_12_4_port, A2 => ab_13_4_port, ZN => 
                           net82635);
   U90 : NAND2_X1 port map( A1 => SUMB_12_5_port, A2 => CARRYB_12_4_port, ZN =>
                           net82633);
   U91 : NAND2_X1 port map( A1 => CARRYB_11_5_port, A2 => SUMB_11_6_port, ZN =>
                           net86250);
   U92 : NAND2_X1 port map( A1 => ab_12_5_port, A2 => CARRYB_11_5_port, ZN => 
                           net86248);
   U93 : NAND2_X1 port map( A1 => CARRYB_10_6_port, A2 => SUMB_10_7_port, ZN =>
                           net86247);
   U94 : NAND2_X1 port map( A1 => ab_11_6_port, A2 => CARRYB_10_6_port, ZN => 
                           net86245);
   U95 : XOR2_X1 port map( A => ab_11_6_port, B => CARRYB_10_6_port, Z => 
                           net86243);
   U96 : NAND2_X1 port map( A1 => CARRYB_9_7_port, A2 => ab_10_7_port, ZN => 
                           net92268);
   U226 : NAND2_X1 port map( A1 => SUMB_9_8_port, A2 => CARRYB_9_7_port, ZN => 
                           net92266);
   U228 : XNOR2_X1 port map( A => net82505, B => SUMB_7_9_port, ZN => 
                           SUMB_8_8_port);
   U231 : XNOR2_X1 port map( A => SUMB_6_10_port, B => net82767, ZN => 
                           SUMB_7_9_port);
   U232 : XNOR2_X1 port map( A => CARRYB_7_8_port, B => ab_8_8_port, ZN => 
                           net82505);
   U233 : CLKBUF_X3 port map( A => net74687, Z => net82987);
   U236 : INV_X1 port map( A => B(7), ZN => net74687);
   U238 : INV_X1 port map( A => B(13), ZN => net74693);
   U239 : INV_X1 port map( A => A(1), ZN => net74665);
   U240 : INV_X1 port map( A => A(2), ZN => net83102);
   U350 : XNOR2_X1 port map( A => ab_0_13_port, B => net82986, ZN => n25);
   U358 : XNOR2_X1 port map( A => CARRYB_6_9_port, B => ab_7_9_port, ZN => 
                           net82767);
   U359 : NAND2_X1 port map( A1 => CARRYB_6_9_port, A2 => ab_7_9_port, ZN => 
                           net82681);
   U360 : NAND2_X1 port map( A1 => SUMB_6_10_port, A2 => CARRYB_6_9_port, ZN =>
                           net82679);
   U361 : NAND2_X1 port map( A1 => CARRYB_5_10_port, A2 => ab_6_10_port, ZN => 
                           net83939);
   U362 : NAND2_X1 port map( A1 => SUMB_5_11_port, A2 => CARRYB_5_10_port, ZN 
                           => net83937);
   U363 : XOR2_X1 port map( A => CARRYB_5_10_port, B => ab_6_10_port, Z => 
                           net83936);
   U364 : XNOR2_X1 port map( A => SUMB_3_12_port, B => net82396, ZN => 
                           SUMB_4_11_port);
   U367 : INV_X1 port map( A => CARRYB_15_1_port, ZN => net82441);
   U368 : XNOR2_X1 port map( A => SUMB_15_1_port, B => net97026, ZN => n41);
   U371 : INV_X1 port map( A => net95080, ZN => net118629);
   U373 : INV_X2 port map( A => net118629, ZN => net118631);
   U375 : XOR2_X1 port map( A => CARRYB_11_7_port, B => ab_12_7_port, Z => n108
                           );
   U376 : XOR2_X1 port map( A => SUMB_11_8_port, B => n108, Z => SUMB_12_7_port
                           );
   U377 : NAND2_X1 port map( A1 => SUMB_11_8_port, A2 => CARRYB_11_7_port, ZN 
                           => n109);
   U378 : NAND2_X1 port map( A1 => SUMB_11_8_port, A2 => ab_12_7_port, ZN => 
                           n110);
   U379 : NAND2_X1 port map( A1 => CARRYB_11_7_port, A2 => ab_12_7_port, ZN => 
                           n111);
   U382 : NOR2_X1 port map( A1 => net74694, A2 => net77075, ZN => n112);
   U383 : INV_X1 port map( A => n112, ZN => n139);
   U384 : XOR2_X1 port map( A => ab_6_14_port, B => ab_5_15_port, Z => n113);
   U385 : XOR2_X1 port map( A => CARRYB_5_14_port, B => n113, Z => 
                           SUMB_6_14_port);
   U386 : NAND2_X1 port map( A1 => CARRYB_5_14_port, A2 => ab_6_14_port, ZN => 
                           n114);
   U387 : NAND2_X1 port map( A1 => CARRYB_5_14_port, A2 => ab_5_15_port, ZN => 
                           n115);
   U388 : NAND2_X1 port map( A1 => ab_6_14_port, A2 => ab_5_15_port, ZN => n116
                           );
   U392 : NOR2_X1 port map( A1 => n187, A2 => net83062, ZN => n117);
   U393 : NOR2_X1 port map( A1 => n141, A2 => TC, ZN => n118);
   U394 : XNOR2_X1 port map( A => SUMB_14_1_port, B => n119, ZN => 
                           SUMB_15_0_port);
   U395 : XNOR2_X1 port map( A => CARRYB_14_0_port, B => ab_15_0_port, ZN => 
                           n119);
   U397 : XOR2_X1 port map( A => CARRYB_9_8_port, B => ab_10_8_port, Z => n120)
                           ;
   U398 : XOR2_X1 port map( A => SUMB_9_9_port, B => n120, Z => SUMB_10_8_port)
                           ;
   U399 : NAND2_X1 port map( A1 => SUMB_9_9_port, A2 => CARRYB_9_8_port, ZN => 
                           n121);
   U400 : NAND2_X1 port map( A1 => SUMB_9_9_port, A2 => ab_10_8_port, ZN => 
                           n122);
   U401 : NAND2_X1 port map( A1 => CARRYB_9_8_port, A2 => ab_10_8_port, ZN => 
                           n123);
   U407 : CLKBUF_X1 port map( A => TC, Z => n125);
   U408 : XOR2_X1 port map( A => ab_3_15_port, B => ab_4_14_port, Z => n126);
   U409 : XOR2_X1 port map( A => CARRYB_3_14_port, B => n126, Z => 
                           SUMB_4_14_port);
   U410 : NAND2_X1 port map( A1 => CARRYB_3_14_port, A2 => ab_3_15_port, ZN => 
                           n127);
   U411 : NAND2_X1 port map( A1 => CARRYB_3_14_port, A2 => ab_4_14_port, ZN => 
                           n128);
   U412 : NAND2_X1 port map( A1 => ab_3_15_port, A2 => ab_4_14_port, ZN => n129
                           );
   U414 : XOR2_X1 port map( A => CARRYB_12_6_port, B => ab_13_6_port, Z => n130
                           );
   U415 : XOR2_X1 port map( A => n130, B => SUMB_12_7_port, Z => SUMB_13_6_port
                           );
   U416 : NAND2_X1 port map( A1 => SUMB_12_7_port, A2 => CARRYB_12_6_port, ZN 
                           => n131);
   U417 : NAND2_X1 port map( A1 => SUMB_12_7_port, A2 => ab_13_6_port, ZN => 
                           n132);
   U418 : NAND2_X1 port map( A1 => CARRYB_12_6_port, A2 => ab_13_6_port, ZN => 
                           n133);
   U422 : NAND2_X1 port map( A1 => SUMB_10_8_port, A2 => CARRYB_10_7_port, ZN 
                           => n135);
   U423 : NAND2_X1 port map( A1 => SUMB_10_8_port, A2 => ab_11_7_port, ZN => 
                           n136);
   U424 : NAND2_X1 port map( A1 => CARRYB_10_7_port, A2 => ab_11_7_port, ZN => 
                           n137);
   U426 : XNOR2_X1 port map( A => n138, B => SUMB_7_10_port, ZN => 
                           SUMB_8_9_port);
   U427 : XNOR2_X1 port map( A => CARRYB_7_9_port, B => ab_8_9_port, ZN => n138
                           );
   U428 : INV_X1 port map( A => B(10), ZN => net82724);
   U429 : INV_X1 port map( A => net77076, ZN => net96980);
   U430 : NAND2_X1 port map( A1 => B(3), A2 => net96980, ZN => n140);
   U431 : INV_X1 port map( A => n140, ZN => ab_1_3_port);
   U432 : INV_X1 port map( A => B(15), ZN => n141);
   U433 : XNOR2_X1 port map( A => CARRYB_2_14_port, B => n142, ZN => 
                           SUMB_3_14_port);
   U434 : XNOR2_X1 port map( A => ab_3_14_port, B => ab_2_15_port, ZN => n142);
   U435 : XNOR2_X1 port map( A => SUMB_3_13_port, B => n143, ZN => 
                           SUMB_4_12_port);
   U436 : XNOR2_X1 port map( A => CARRYB_3_12_port, B => ab_4_12_port, ZN => 
                           n143);
   U437 : XOR2_X1 port map( A => CARRYB_13_5_port, B => ab_14_5_port, Z => n144
                           );
   U438 : XOR2_X1 port map( A => SUMB_13_6_port, B => n144, Z => SUMB_14_5_port
                           );
   U439 : NAND2_X1 port map( A1 => SUMB_13_6_port, A2 => CARRYB_13_5_port, ZN 
                           => n145);
   U440 : NAND2_X1 port map( A1 => SUMB_13_6_port, A2 => ab_14_5_port, ZN => 
                           n146);
   U441 : NAND2_X1 port map( A1 => CARRYB_13_5_port, A2 => ab_14_5_port, ZN => 
                           n147);
   U445 : NAND2_X1 port map( A1 => SUMB_14_5_port, A2 => CARRYB_14_4_port, ZN 
                           => n149);
   U446 : NAND2_X1 port map( A1 => SUMB_14_5_port, A2 => ab_15_4_port, ZN => 
                           n150);
   U447 : NAND2_X1 port map( A1 => CARRYB_14_4_port, A2 => ab_15_4_port, ZN => 
                           n151);
   U449 : XNOR2_X1 port map( A => CARRYB_14_3_port, B => ab_15_3_port, ZN => 
                           n152);
   U454 : CLKBUF_X1 port map( A => net74665, Z => net77076);
   U455 : NAND2_X1 port map( A1 => SUMB_7_10_port, A2 => CARRYB_7_9_port, ZN =>
                           n153);
   U456 : NAND2_X1 port map( A1 => SUMB_7_10_port, A2 => ab_8_9_port, ZN => 
                           n154);
   U457 : NAND2_X1 port map( A1 => CARRYB_7_9_port, A2 => ab_8_9_port, ZN => 
                           n155);
   U459 : XOR2_X1 port map( A => CARRYB_11_6_port, B => ab_12_6_port, Z => n156
                           );
   U460 : XOR2_X1 port map( A => n156, B => SUMB_11_7_port, Z => SUMB_12_6_port
                           );
   U461 : NAND2_X1 port map( A1 => SUMB_11_7_port, A2 => CARRYB_11_6_port, ZN 
                           => n157);
   U462 : NAND2_X1 port map( A1 => SUMB_11_7_port, A2 => ab_12_6_port, ZN => 
                           n158);
   U463 : NAND2_X1 port map( A1 => CARRYB_11_6_port, A2 => ab_12_6_port, ZN => 
                           n159);
   U465 : INV_X1 port map( A => CARRYB_15_4_port, ZN => n168);
   U467 : NAND2_X1 port map( A1 => CARRYB_3_12_port, A2 => SUMB_3_13_port, ZN 
                           => n161);
   U468 : NAND2_X1 port map( A1 => SUMB_3_13_port, A2 => ab_4_12_port, ZN => 
                           n162);
   U469 : NAND2_X1 port map( A1 => CARRYB_3_12_port, A2 => ab_4_12_port, ZN => 
                           n163);
   U472 : XNOR2_X1 port map( A => SUMB_14_4_port, B => n152, ZN => 
                           SUMB_15_3_port);
   U473 : INV_X1 port map( A => CARRYB_15_3_port, ZN => n166);
   U475 : XNOR2_X1 port map( A => n166, B => SUMB_15_4_port, ZN => n35);
   U477 : NAND2_X1 port map( A1 => SUMB_9_8_port, A2 => ab_10_7_port, ZN => 
                           n167);
   U479 : XNOR2_X1 port map( A => SUMB_15_5_port, B => n168, ZN => n50);
   U480 : NAND2_X1 port map( A1 => SUMB_14_1_port, A2 => CARRYB_14_0_port, ZN 
                           => net88955);
   U481 : NAND2_X1 port map( A1 => SUMB_14_1_port, A2 => ab_15_0_port, ZN => 
                           net88956);
   U482 : NAND2_X1 port map( A1 => CARRYB_14_0_port, A2 => ab_15_0_port, ZN => 
                           net88957);
   U487 : NAND2_X1 port map( A1 => SUMB_14_4_port, A2 => CARRYB_14_3_port, ZN 
                           => n170);
   U488 : NAND2_X1 port map( A1 => SUMB_14_4_port, A2 => ab_15_3_port, ZN => 
                           n171);
   U489 : NAND2_X1 port map( A1 => CARRYB_14_3_port, A2 => ab_15_3_port, ZN => 
                           n172);
   U491 : XNOR2_X1 port map( A => n173, B => n17, ZN => SUMB_2_14_port);
   U492 : XNOR2_X1 port map( A => ab_1_15_port, B => ab_2_14_port, ZN => n173);
   U494 : XOR2_X1 port map( A => net86243, B => SUMB_10_7_port, Z => 
                           SUMB_11_6_port);
   U495 : NAND2_X1 port map( A1 => ab_11_6_port, A2 => SUMB_10_7_port, ZN => 
                           n174);
   U497 : NAND2_X1 port map( A1 => ab_12_5_port, A2 => SUMB_11_6_port, ZN => 
                           n175);
   U499 : XOR2_X1 port map( A => SUMB_5_11_port, B => net83936, Z => 
                           SUMB_6_10_port);
   U500 : NAND2_X1 port map( A1 => SUMB_5_11_port, A2 => ab_6_10_port, ZN => 
                           n176);
   U502 : NOR2_X1 port map( A1 => n177, A2 => n243, ZN => n8);
   U503 : NAND2_X1 port map( A1 => n185, A2 => net83064, ZN => n177);
   U511 : CLKBUF_X3 port map( A => n243, Z => n184);
   U513 : INV_X1 port map( A => n185, ZN => n223);
   U514 : CLKBUF_X1 port map( A => net82475, Z => net83064);
   U515 : CLKBUF_X1 port map( A => net77069, Z => net83062);
   U516 : CLKBUF_X3 port map( A => n276, Z => n186);
   U517 : INV_X1 port map( A => B(5), ZN => n276);
   U518 : XNOR2_X1 port map( A => n223, B => ab_0_9_port, ZN => n22);
   U520 : INV_X1 port map( A => B(4), ZN => n187);
   U522 : XNOR2_X1 port map( A => net82980, B => ab_1_10_port, ZN => n21);
   U524 : XNOR2_X1 port map( A => n140, B => n117, ZN => n18);
   U525 : CLKBUF_X3 port map( A => n275, Z => n189);
   U526 : INV_X1 port map( A => B(6), ZN => n275);
   U530 : CLKBUF_X1 port map( A => n274, Z => n192);
   U531 : INV_X1 port map( A => B(8), ZN => n274);
   U534 : XNOR2_X1 port map( A => n194, B => n232, ZN => SUMB_2_13_port);
   U535 : XOR2_X1 port map( A => n245, B => n139, Z => n194);
   U536 : INV_X1 port map( A => A(3), ZN => net82975);
   U537 : INV_X1 port map( A => A(3), ZN => net82976);
   U541 : XNOR2_X1 port map( A => net82942, B => SUMB_15_3_port, ZN => n49);
   U543 : XNOR2_X1 port map( A => n293, B => n197, ZN => SUMB_2_9_port);
   U544 : XNOR2_X1 port map( A => n10, B => ab_2_9_port, ZN => n197);
   U545 : XOR2_X1 port map( A => CARRYB_13_0_port, B => ab_14_0_port, Z => n198
                           );
   U546 : XOR2_X1 port map( A => SUMB_13_1_port, B => n198, Z => A1_12_port);
   U547 : NAND2_X1 port map( A1 => SUMB_13_1_port, A2 => CARRYB_13_0_port, ZN 
                           => n199);
   U548 : NAND2_X1 port map( A1 => SUMB_13_1_port, A2 => ab_14_0_port, ZN => 
                           n200);
   U549 : NAND2_X1 port map( A1 => CARRYB_13_0_port, A2 => ab_14_0_port, ZN => 
                           n201);
   U552 : XNOR2_X1 port map( A => n245, B => n139, ZN => n204);
   U553 : XNOR2_X1 port map( A => SUMB_12_5_port, B => net82778, ZN => net82876
                           );
   U554 : NAND2_X1 port map( A1 => n21, A2 => n10, ZN => n205);
   U555 : NAND2_X1 port map( A1 => n293, A2 => ab_2_9_port, ZN => n206);
   U556 : NAND2_X1 port map( A1 => n10, A2 => n297, ZN => n207);
   U558 : NAND2_X1 port map( A1 => n17, A2 => ab_1_15_port, ZN => n208);
   U559 : NAND2_X1 port map( A1 => n17, A2 => ab_2_14_port, ZN => n209);
   U560 : NAND2_X1 port map( A1 => ab_1_15_port, A2 => ab_2_14_port, ZN => n210
                           );
   U563 : INV_X1 port map( A => B(0), ZN => net74680);
   U565 : XNOR2_X1 port map( A => n211, B => ab_1_9_port, ZN => n24);
   U566 : OR2_X1 port map( A1 => net77069, A2 => net74690, ZN => n211);
   U567 : XNOR2_X1 port map( A => n27, B => n212, ZN => SUMB_2_6_port);
   U568 : XNOR2_X1 port map( A => n14, B => ab_2_6_port, ZN => n212);
   U569 : NAND2_X1 port map( A1 => n27, A2 => n14, ZN => n213);
   U570 : NAND2_X1 port map( A1 => n27, A2 => ab_2_6_port, ZN => n214);
   U571 : NAND2_X1 port map( A1 => n14, A2 => ab_2_6_port, ZN => n215);
   U574 : INV_X1 port map( A => B(10), ZN => net74690);
   U576 : NAND2_X1 port map( A1 => SUMB_6_10_port, A2 => ab_7_9_port, ZN => 
                           n218);
   U578 : INV_X1 port map( A => net74665, ZN => net82622);
   U579 : NAND2_X1 port map( A1 => CARRYB_2_14_port, A2 => ab_3_14_port, ZN => 
                           n219);
   U580 : NAND2_X1 port map( A1 => CARRYB_2_14_port, A2 => ab_2_15_port, ZN => 
                           n220);
   U581 : NAND2_X1 port map( A1 => ab_3_14_port, A2 => ab_2_15_port, ZN => n221
                           );
   U583 : NAND2_X1 port map( A1 => SUMB_12_5_port, A2 => ab_13_4_port, ZN => 
                           n222);
   U586 : INV_X1 port map( A => net74664, ZN => net82475);
   U587 : XNOR2_X1 port map( A => net82876, B => net82608, ZN => SUMB_14_3_port
                           );
   U588 : NAND2_X1 port map( A1 => net82876, A2 => ab_14_3_port, ZN => n224);
   U590 : XNOR2_X1 port map( A => n245, B => n139, ZN => n31);
   U591 : XOR2_X1 port map( A => n267, B => net118631, Z => n225);
   U592 : XOR2_X1 port map( A => SUMB_15_0_port, B => n225, Z => A1_13_port);
   U593 : NAND2_X1 port map( A1 => SUMB_15_0_port, A2 => n267, ZN => n226);
   U594 : NAND2_X1 port map( A1 => SUMB_15_0_port, A2 => net118631, ZN => n227)
                           ;
   U595 : NAND2_X1 port map( A1 => n267, A2 => net118631, ZN => n228);
   U597 : CLKBUF_X1 port map( A => net74694, Z => net82535);
   U598 : NAND2_X1 port map( A1 => SUMB_7_9_port, A2 => CARRYB_7_8_port, ZN => 
                           n229);
   U599 : NAND2_X1 port map( A1 => SUMB_7_9_port, A2 => ab_8_8_port, ZN => n230
                           );
   U600 : NAND2_X1 port map( A1 => CARRYB_7_8_port, A2 => ab_8_8_port, ZN => 
                           n231);
   U602 : XOR2_X1 port map( A => n12, B => ab_2_13_port, Z => n232);
   U603 : NAND2_X1 port map( A1 => n31, A2 => n12, ZN => n233);
   U604 : NAND2_X1 port map( A1 => n204, A2 => ab_2_13_port, ZN => n234);
   U605 : NAND2_X1 port map( A1 => n12, A2 => ab_2_13_port, ZN => n235);
   U609 : XNOR2_X1 port map( A => SUMB_15_2_port, B => net82441, ZN => n34);
   U610 : NOR2_X1 port map( A1 => net74693, A2 => net77075, ZN => n238);
   U612 : XNOR2_X1 port map( A => SUMB_2_13_port, B => net82414, ZN => 
                           SUMB_3_12_port);
   U613 : NAND2_X1 port map( A1 => ab_3_12_port, A2 => SUMB_2_13_port, ZN => 
                           n239);
   U615 : NAND2_X1 port map( A1 => ab_4_11_port, A2 => CARRYB_3_11_port, ZN => 
                           n240);
   U616 : NAND2_X1 port map( A1 => ab_4_11_port, A2 => SUMB_3_12_port, ZN => 
                           n241);
   U617 : NAND2_X1 port map( A1 => CARRYB_3_11_port, A2 => SUMB_3_12_port, ZN 
                           => n242);
   U619 : CLKBUF_X3 port map( A => net74664, Z => net77069);
   U620 : NOR2_X1 port map( A1 => n272, A2 => n125, ZN => net82309);
   U621 : INV_X2 port map( A => B(3), ZN => n278);
   U622 : INV_X2 port map( A => A(4), ZN => n290);
   U623 : INV_X1 port map( A => B(9), ZN => n243);
   U631 : CLKBUF_X1 port map( A => n289, Z => n265);
   U632 : CLKBUF_X1 port map( A => n289, Z => n266);
   U643 : CLKBUF_X1 port map( A => ZA, Z => n267);
   U655 : INV_X1 port map( A => A(15), ZN => n281);
   U656 : INV_X1 port map( A => A(6), ZN => n289);
   U657 : INV_X1 port map( A => A(10), ZN => n286);
   U658 : INV_X1 port map( A => A(5), ZN => net74669);
   U659 : INV_X1 port map( A => A(9), ZN => net74673);
   U660 : INV_X1 port map( A => A(8), ZN => n287);
   U661 : INV_X1 port map( A => A(11), ZN => n285);
   U662 : INV_X1 port map( A => A(14), ZN => n282);
   U663 : INV_X1 port map( A => A(7), ZN => n288);
   U665 : INV_X1 port map( A => A(13), ZN => n283);
   U666 : INV_X1 port map( A => A(12), ZN => n284);
   U667 : CLKBUF_X1 port map( A => net82309, Z => net76791);
   U668 : MUX2_X2 port map( A => n98, B => net95080, S => net77069, Z => n245);
   U669 : INV_X1 port map( A => B(15), ZN => n272);
   U670 : INV_X1 port map( A => n125, ZN => n291);
   FS_1 : ALU_N32_DW01_add_0 port map( A(29) => n63, A(28) => n62, A(27) => n40
                           , A(26) => n54, A(25) => n39, A(24) => n53, A(23) =>
                           n38, A(22) => n52, A(21) => n37, A(20) => n51, A(19)
                           => n36, A(18) => n50, A(17) => n35, A(16) => n49, 
                           A(15) => n34, A(14) => n41, A(13) => A1_13_port, 
                           A(12) => A1_12_port, A(11) => A1_11_port, A(10) => 
                           A1_10_port, A(9) => A1_9_port, A(8) => A1_8_port, 
                           A(7) => A1_7_port, A(6) => A1_6_port, A(5) => 
                           A1_5_port, A(4) => A1_4_port, A(3) => A1_3_port, 
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(29) => n32, B(28) => n61, B(27) => n48,
                           B(26) => n60, B(25) => n47, B(24) => n59, B(23) => 
                           n46, B(22) => n58, B(21) => n45, B(20) => n57, B(19)
                           => n44, B(18) => n56, B(17) => n43, B(16) => n55, 
                           B(15) => n42, B(14) => A2_14_port, B(13) => n101, 
                           B(12) => n101, B(11) => n101, B(10) => n101, B(9) =>
                           n101, B(8) => n101, B(7) => n101, B(6) => n101, B(5)
                           => n101, B(4) => n101, B(3) => n101, B(2) => n101, 
                           B(1) => n101, B(0) => n100, CI => n100, SUM(29) => 
                           PRODUCT(31), SUM(28) => PRODUCT(30), SUM(27) => 
                           PRODUCT(29), SUM(26) => PRODUCT(28), SUM(25) => 
                           PRODUCT(27), SUM(24) => PRODUCT(26), SUM(23) => 
                           PRODUCT(25), SUM(22) => PRODUCT(24), SUM(21) => 
                           PRODUCT(23), SUM(20) => PRODUCT(22), SUM(19) => 
                           PRODUCT(21), SUM(18) => PRODUCT(20), SUM(17) => 
                           PRODUCT(19), SUM(16) => PRODUCT(18), SUM(15) => 
                           PRODUCT(17), SUM(14) => PRODUCT(16), SUM(13) => 
                           PRODUCT(15), SUM(12) => PRODUCT(14), SUM(11) => 
                           PRODUCT(13), SUM(10) => PRODUCT(12), SUM(9) => 
                           PRODUCT(11), SUM(8) => PRODUCT(10), SUM(7) => 
                           PRODUCT(9), SUM(6) => PRODUCT(8), SUM(5) => 
                           PRODUCT(7), SUM(4) => PRODUCT(6), SUM(3) => 
                           PRODUCT(5), SUM(2) => PRODUCT(4), SUM(1) => 
                           PRODUCT(3), SUM(0) => PRODUCT(2), CO => n_1020);
   U2 : AND2_X1 port map( A1 => ab_1_9_port, A2 => ab_0_10_port, ZN => n10);
   U3 : INV_X2 port map( A => B(1), ZN => n280);
   U4 : MUX2_X1 port map( A => net76791, B => net118631, S => net82975, Z => 
                           ab_3_15_port);
   U5 : MUX2_X1 port map( A => net82309, B => net95080, S => net83102, Z => 
                           ab_2_15_port);
   U6 : NAND3_X1 port map( A1 => n153, A2 => n154, A3 => n155, ZN => 
                           CARRYB_8_9_port);
   U7 : CLKBUF_X1 port map( A => net74693, Z => net118627);
   U8 : AND2_X1 port map( A1 => TC, A2 => B(15), ZN => net95080);
   U9 : AND2_X1 port map( A1 => CARRYB_15_4_port, A2 => SUMB_15_5_port, ZN => 
                           n44);
   U10 : CLKBUF_X1 port map( A => net74665, Z => net77075);
   U11 : AND2_X1 port map( A1 => B(4), A2 => net96980, ZN => n292);
   U12 : MUX2_X1 port map( A => n118, B => net95080, S => net77075, Z => 
                           ab_1_15_port);
   U13 : AND2_X1 port map( A1 => net82475, A2 => B(12), ZN => ab_0_12_port);
   U14 : XNOR2_X1 port map( A => net82980, B => ab_1_10_port, ZN => n293);
   U15 : BUF_X1 port map( A => A(0), Z => net83044);
   U16 : XNOR2_X1 port map( A => SUMB_9_8_port, B => n294, ZN => SUMB_10_7_port
                           );
   U17 : XNOR2_X1 port map( A => CARRYB_9_7_port, B => ab_10_7_port, ZN => n294
                           );
   U20 : XNOR2_X1 port map( A => SUMB_14_5_port, B => n295, ZN => 
                           SUMB_15_4_port);
   U21 : XNOR2_X1 port map( A => CARRYB_14_4_port, B => ab_15_4_port, ZN => 
                           n295);
   U22 : XNOR2_X1 port map( A => n296, B => ab_0_7_port, ZN => n28);
   U25 : OR2_X1 port map( A1 => n275, A2 => net77076, ZN => n296);
   U27 : BUF_X1 port map( A => A(1), Z => n102);
   U30 : NOR2_X1 port map( A1 => n243, A2 => net83102, ZN => n297);
   U31 : XNOR2_X1 port map( A => SUMB_10_8_port, B => n298, ZN => 
                           SUMB_11_7_port);
   U33 : XNOR2_X1 port map( A => CARRYB_10_7_port, B => ab_11_7_port, ZN => 
                           n298);
   U36 : XNOR2_X1 port map( A => n299, B => SUMB_14_6_port, ZN => 
                           SUMB_15_5_port);
   U42 : XNOR2_X1 port map( A => ab_15_5_port, B => CARRYB_14_5_port, ZN => 
                           n299);
   U43 : AND2_X1 port map( A1 => net82534, A2 => n238, ZN => n12);
   U44 : XOR2_X1 port map( A => ab_1_11_port, B => ab_0_12_port, Z => n23);
   U45 : XOR2_X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, Z => n300)
                           ;
   U46 : XOR2_X1 port map( A => n300, B => SUMB_13_7_port, Z => SUMB_14_6_port)
                           ;
   U47 : NAND2_X1 port map( A1 => ab_14_6_port, A2 => CARRYB_13_6_port, ZN => 
                           n301);
   U48 : NAND2_X1 port map( A1 => ab_14_6_port, A2 => SUMB_13_7_port, ZN => 
                           n302);
   U49 : NAND2_X1 port map( A1 => CARRYB_13_6_port, A2 => SUMB_13_7_port, ZN =>
                           n303);
   U56 : NAND3_X1 port map( A1 => n301, A2 => n302, A3 => n303, ZN => 
                           CARRYB_14_6_port);
   U57 : NAND2_X1 port map( A1 => ab_15_5_port, A2 => CARRYB_14_5_port, ZN => 
                           n304);
   U58 : NAND2_X1 port map( A1 => ab_15_5_port, A2 => SUMB_14_6_port, ZN => 
                           n305);
   U59 : NAND2_X1 port map( A1 => CARRYB_14_5_port, A2 => SUMB_14_6_port, ZN =>
                           n306);
   U60 : NAND3_X1 port map( A1 => n304, A2 => n305, A3 => n306, ZN => 
                           CARRYB_15_5_port);
   U61 : INV_X2 port map( A => net82651, ZN => net82653);
   U62 : INV_X1 port map( A => CARRYB_15_2_port, ZN => net82942);
   U66 : AND2_X1 port map( A1 => n245, A2 => n112, ZN => n17);
   U73 : AND2_X1 port map( A1 => n102, A2 => B(11), ZN => ab_1_11_port);
   U74 : NAND3_X1 port map( A1 => net82385, A2 => n239, A3 => net82387, ZN => 
                           CARRYB_3_12_port);
   U75 : MUX2_X1 port map( A => net76791, B => net118631, S => n289, Z => 
                           ab_6_15_port);
   U77 : NAND3_X1 port map( A1 => n114, A2 => n115, A3 => n116, ZN => 
                           CARRYB_6_14_port);
   U80 : NAND3_X1 port map( A1 => n229, A2 => n230, A3 => n231, ZN => 
                           CARRYB_8_8_port);
   U81 : MUX2_X1 port map( A => net76791, B => net118631, S => net74673, Z => 
                           ab_9_15_port);
   U107 : NAND3_X1 port map( A1 => n131, A2 => n132, A3 => n133, ZN => 
                           CARRYB_13_6_port);
   U123 : NAND3_X1 port map( A1 => net86248, A2 => n175, A3 => net86250, ZN => 
                           CARRYB_12_5_port);
   U139 : MUX2_X1 port map( A => net76791, B => net118631, S => n284, Z => 
                           ab_12_15_port);
   U155 : MUX2_X1 port map( A => n99, B => ZA, S => n181, Z => ab_15_2_port);
   U171 : NAND3_X1 port map( A1 => n149, A2 => n150, A3 => n151, ZN => 
                           CARRYB_15_4_port);
   U187 : AND2_X1 port map( A1 => CARRYB_15_13_port, A2 => SUMB_15_14_port, ZN 
                           => n61);
   U203 : AND2_X1 port map( A1 => CARRYB_15_2_port, A2 => SUMB_15_3_port, ZN =>
                           n43);
   U219 : AND2_X1 port map( A1 => CARRYB_15_8_port, A2 => SUMB_15_9_port, ZN =>
                           n46);
   U227 : AND2_X1 port map( A1 => CARRYB_15_9_port, A2 => SUMB_15_10_port, ZN 
                           => n59);
   U235 : NAND3_X1 port map( A1 => n219, A2 => n220, A3 => n221, ZN => 
                           CARRYB_3_14_port);
   U237 : AND2_X1 port map( A1 => B(14), A2 => net83044, ZN => net82534);
   U242 : AND2_X1 port map( A1 => B(13), A2 => net83044, ZN => ab_0_13_port);
   U243 : AND2_X1 port map( A1 => A(1), A2 => B(12), ZN => ab_1_12_port);
   U244 : NAND3_X1 port map( A1 => n234, A2 => n233, A3 => n235, ZN => 
                           CARRYB_2_13_port);
   U245 : AND2_X1 port map( A1 => ab_0_11_port, A2 => ab_1_10_port, ZN => n7);
   U246 : AND2_X1 port map( A1 => net82622, A2 => B(9), ZN => ab_1_9_port);
   U247 : NAND3_X1 port map( A1 => n240, A2 => n241, A3 => n242, ZN => 
                           CARRYB_4_11_port);
   U248 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n14);
   U249 : AND2_X1 port map( A1 => ab_0_8_port, A2 => ab_1_7_port, ZN => n13);
   U250 : MUX2_X1 port map( A => net82309, B => net118631, S => n287, Z => 
                           ab_8_15_port);
   U252 : NAND3_X1 port map( A1 => net86245, A2 => n174, A3 => net86247, ZN => 
                           CARRYB_11_6_port);
   U253 : NAND3_X1 port map( A1 => net92266, A2 => n167, A3 => net92268, ZN => 
                           CARRYB_10_7_port);
   U254 : NAND3_X1 port map( A1 => n170, A2 => n171, A3 => n172, ZN => 
                           CARRYB_15_3_port);
   U255 : MUX2_X1 port map( A => net76791, B => net118631, S => n285, Z => 
                           ab_11_15_port);
   U256 : MUX2_X1 port map( A => n99, B => ZA, S => n280, Z => ab_15_1_port);
   U257 : NAND3_X1 port map( A1 => n109, A2 => n110, A3 => n111, ZN => 
                           CARRYB_12_7_port);
   U268 : AND2_X1 port map( A1 => B(2), A2 => net96980, ZN => ab_1_2_port);
   U284 : NAND3_X1 port map( A1 => n199, A2 => n200, A3 => n201, ZN => 
                           CARRYB_14_0_port);
   U300 : MUX2_X1 port map( A => n99, B => ZA, S => n186, Z => ab_15_5_port);
   U316 : NAND3_X1 port map( A1 => n145, A2 => n146, A3 => n147, ZN => 
                           CARRYB_14_5_port);
   U332 : AND2_X1 port map( A1 => CARRYB_15_7_port, A2 => SUMB_15_8_port, ZN =>
                           n58);
   U348 : MUX2_X1 port map( A => n99, B => n267, S => net82724, Z => 
                           ab_15_10_port);
   U351 : MUX2_X1 port map( A => n99, B => ZA, S => net82653, Z => 
                           ab_15_11_port);
   U352 : MUX2_X1 port map( A => net76791, B => net118631, S => n282, Z => 
                           ab_14_15_port);
   U365 : MUX2_X1 port map( A => n99, B => ZA, S => net82535, Z => 
                           ab_15_14_port);
   U366 : MUX2_X1 port map( A => n99, B => ZA, S => net97008, Z => 
                           ab_15_12_port);
   U369 : MUX2_X1 port map( A => n99, B => ZA, S => net118627, Z => 
                           ab_15_13_port);
   U370 : AND2_X1 port map( A1 => CARRYB_15_11_port, A2 => SUMB_15_12_port, ZN 
                           => n60);
   U372 : AND2_X1 port map( A1 => CARRYB_15_14_port, A2 => SUMB_15_15_port, ZN 
                           => n32);
   U374 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n4);
   U380 : AND2_X1 port map( A1 => n102, A2 => B(10), ZN => ab_1_10_port);
   U381 : NAND3_X1 port map( A1 => n208, A2 => n209, A3 => n210, ZN => 
                           CARRYB_2_14_port);
   U389 : AND2_X1 port map( A1 => ab_1_11_port, A2 => ab_0_12_port, ZN => n9);
   U390 : AND2_X1 port map( A1 => ab_1_12_port, A2 => ab_0_13_port, ZN => n11);
   U391 : MUX2_X1 port map( A => net82309, B => net118631, S => net74669, Z => 
                           ab_5_15_port);
   U396 : MUX2_X1 port map( A => net76791, B => net118631, S => n290, Z => 
                           ab_4_15_port);
   U402 : NAND3_X1 port map( A1 => n127, A2 => n128, A3 => n129, ZN => 
                           CARRYB_4_14_port);
   U403 : AND2_X1 port map( A1 => net82622, A2 => B(8), ZN => n185);
   U404 : NAND3_X1 port map( A1 => n206, A2 => n205, A3 => n207, ZN => 
                           CARRYB_2_9_port);
   U405 : NAND3_X1 port map( A1 => n161, A2 => n162, A3 => n163, ZN => 
                           CARRYB_4_12_port);
   U406 : MUX2_X1 port map( A => net76791, B => net118631, S => n288, Z => 
                           ab_7_15_port);
   U413 : AND2_X1 port map( A1 => B(7), A2 => net82622, ZN => ab_1_7_port);
   U419 : NAND3_X1 port map( A1 => net82679, A2 => n218, A3 => net82681, ZN => 
                           CARRYB_7_9_port);
   U420 : NAND3_X1 port map( A1 => n176, A2 => net83937, A3 => net83939, ZN => 
                           CARRYB_6_10_port);
   U421 : NAND3_X1 port map( A1 => n214, A2 => n213, A3 => n215, ZN => 
                           CARRYB_2_6_port);
   U425 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n15);
   U442 : NAND3_X1 port map( A1 => n121, A2 => n122, A3 => n123, ZN => 
                           CARRYB_10_8_port);
   U443 : MUX2_X1 port map( A => net82309, B => net118631, S => n286, Z => 
                           ab_10_15_port);
   U444 : AND2_X1 port map( A1 => ab_0_5_port, A2 => n292, ZN => n16);
   U448 : NAND3_X1 port map( A1 => n135, A2 => n136, A3 => n137, ZN => 
                           CARRYB_11_7_port);
   U450 : NAND3_X1 port map( A1 => n157, A2 => n158, A3 => n159, ZN => 
                           CARRYB_12_6_port);
   U451 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n3);
   U452 : AND2_X1 port map( A1 => CARRYB_15_1_port, A2 => SUMB_15_2_port, ZN =>
                           n55);
   U453 : NAND3_X1 port map( A1 => net82595, A2 => n224, A3 => net82597, ZN => 
                           CARRYB_14_3_port);
   U458 : MUX2_X1 port map( A => n99, B => ZA, S => n278, Z => ab_15_3_port);
   U464 : AND2_X1 port map( A1 => SUMB_15_4_port, A2 => CARRYB_15_3_port, ZN =>
                           n56);
   U466 : MUX2_X1 port map( A => n99, B => ZA, S => n248, Z => ab_15_4_port);
   U470 : NAND3_X1 port map( A1 => net82633, A2 => n222, A3 => net82635, ZN => 
                           CARRYB_13_4_port);
   U471 : MUX2_X1 port map( A => n99, B => ZA, S => net74680, Z => ab_15_0_port
                           );
   U474 : AND3_X1 port map( A1 => net88955, A2 => net88956, A3 => net88957, ZN 
                           => net97026);
   U476 : AND2_X1 port map( A1 => SUMB_15_1_port, A2 => CARRYB_15_0_port, ZN =>
                           n42);
   U478 : NAND3_X1 port map( A1 => net88956, A2 => net88955, A3 => net88957, ZN
                           => CARRYB_15_0_port);
   U483 : MUX2_X1 port map( A => n99, B => ZA, S => n189, Z => ab_15_6_port);
   U484 : MUX2_X1 port map( A => n99, B => n267, S => n184, Z => ab_15_9_port);
   U485 : MUX2_X1 port map( A => net82309, B => net118631, S => n283, Z => 
                           ab_13_15_port);
   U486 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U490 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U493 : NAND3_X1 port map( A1 => n226, A2 => n227, A3 => n228, ZN => 
                           A2_14_port);
   U496 : MUX2_X1 port map( A => n99, B => n267, S => n192, Z => ab_15_8_port);
   U498 : MUX2_X1 port map( A => n99, B => n267, S => net82987, Z => 
                           ab_15_7_port);
   U501 : AND2_X1 port map( A1 => CARRYB_15_6_port, A2 => SUMB_15_7_port, ZN =>
                           n45);
   U504 : AND2_X1 port map( A1 => CARRYB_15_5_port, A2 => SUMB_15_6_port, ZN =>
                           n57);
   U505 : AND2_X1 port map( A1 => CARRYB_15_10_port, A2 => SUMB_15_11_port, ZN 
                           => n47);
   U506 : AND2_X1 port map( A1 => CARRYB_15_12_port, A2 => SUMB_15_13_port, ZN 
                           => n48);
   U507 : INV_X2 port map( A => B(2), ZN => n181);
   U508 : CLKBUF_X3 port map( A => n187, Z => n248);

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_cmp6_1 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end ALU_N32_DW01_cmp6_1;

architecture SYN_rpl of ALU_N32_DW01_cmp6_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n202, GE_port, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n161, n162, n163, n164, 
      n167, n168, n169, n170, n173, n174, n175, n176, n179, n180, n181, n182, 
      n185, n186, n187, n188, n191, n192, n193, n194, n197, n198, n200, n201, 
      n199, n196, n195, n190, n189, n184, n183, n178, n177, n172, n171, n166, 
      n165, n160, LE_port, n204, n205, n206, n207, n208, n209, n210, n211, n212
      , n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265 : std_logic;

begin
   LE <= LE_port;
   GE <= GE_port;
   
   U65 : AOI21_X1 port map( B1 => n65, B2 => n205, A => n66, ZN => GE_port);
   U66 : AOI22_X1 port map( A1 => B(30), A2 => n236, B1 => n68, B2 => n69, ZN 
                           => n67);
   U67 : AOI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n68);
   U68 : AOI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n70);
   U69 : AOI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n73);
   U70 : AOI21_X1 port map( B1 => n79, B2 => n209, A => n210, ZN => n76);
   U71 : AOI21_X1 port map( B1 => n82, B2 => n83, A => n84, ZN => n79);
   U72 : AOI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n82);
   U73 : AOI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n85);
   U74 : AOI21_X1 port map( B1 => n91, B2 => n213, A => n214, ZN => n88);
   U75 : AOI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n91);
   U76 : AOI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n94);
   U77 : AOI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n97);
   U78 : AOI21_X1 port map( B1 => n103, B2 => n217, A => n218, ZN => n100);
   U79 : AOI21_X1 port map( B1 => n106, B2 => n107, A => n108, ZN => n103);
   U80 : AOI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n106);
   U81 : AOI21_X1 port map( B1 => n112, B2 => n113, A => n114, ZN => n109);
   U82 : AOI21_X1 port map( B1 => n115, B2 => n221, A => n222, ZN => n112);
   U83 : AOI21_X1 port map( B1 => n118, B2 => n119, A => n120, ZN => n115);
   U84 : AOI21_X1 port map( B1 => n121, B2 => n122, A => n123, ZN => n118);
   U85 : AOI21_X1 port map( B1 => n124, B2 => n125, A => n126, ZN => n121);
   U86 : AOI21_X1 port map( B1 => n127, B2 => n225, A => n226, ZN => n124);
   U87 : AOI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => n127);
   U88 : AOI21_X1 port map( B1 => n133, B2 => n134, A => n135, ZN => n130);
   U89 : AOI21_X1 port map( B1 => n136, B2 => n137, A => n138, ZN => n133);
   U90 : AOI21_X1 port map( B1 => n139, B2 => n229, A => n230, ZN => n136);
   U91 : AOI21_X1 port map( B1 => n142, B2 => n143, A => n144, ZN => n139);
   U92 : AOI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n142);
   U93 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U94 : AOI21_X1 port map( B1 => n151, B2 => n152, A => n233, ZN => n148);
   U95 : AOI22_X1 port map( A1 => n154, A2 => n235, B1 => A(1), B2 => n155, ZN 
                           => n151);
   U96 : OR2_X1 port map( A1 => n155, A2 => A(1), ZN => n154);
   U97 : NAND2_X1 port map( A1 => B(0), A2 => n265, ZN => n155);
   U98 : OAI21_X1 port map( B1 => n66, B2 => n156, A => n65, ZN => n202);
   U99 : NAND2_X1 port map( A1 => A(31), A2 => n204, ZN => n65);
   U100 : AOI22_X1 port map( A1 => A(30), A2 => n206, B1 => n157, B2 => n69, ZN
                           => n156);
   U101 : XOR2_X1 port map( A => A(30), B => n206, Z => n69);
   U102 : AOI21_X1 port map( B1 => n158, B2 => n159, A => n207, ZN => n157);
   U103 : NAND2_X1 port map( A1 => B(29), A2 => n237, ZN => n71);
   U105 : NOR2_X1 port map( A1 => n162, A2 => n75, ZN => n74);
   U107 : NAND2_X1 port map( A1 => B(27), A2 => n239, ZN => n77);
   U108 : NAND2_X1 port map( A1 => n208, A2 => n163, ZN => n161);
   U109 : NOR2_X1 port map( A1 => n239, A2 => B(27), ZN => n78);
   U111 : NAND2_X1 port map( A1 => B(25), A2 => n241, ZN => n83);
   U112 : NAND2_X1 port map( A1 => n163, A2 => n80, ZN => n81);
   U113 : NAND2_X1 port map( A1 => B(26), A2 => n240, ZN => n80);
   U114 : OR2_X1 port map( A1 => n240, A2 => B(26), ZN => n163);
   U116 : NOR2_X1 port map( A1 => n168, A2 => n87, ZN => n86);
   U118 : NAND2_X1 port map( A1 => B(23), A2 => n243, ZN => n89);
   U119 : NAND2_X1 port map( A1 => n212, A2 => n169, ZN => n167);
   U120 : NOR2_X1 port map( A1 => n243, A2 => B(23), ZN => n90);
   U122 : NAND2_X1 port map( A1 => B(21), A2 => n245, ZN => n95);
   U123 : NAND2_X1 port map( A1 => n169, A2 => n92, ZN => n93);
   U124 : NAND2_X1 port map( A1 => B(22), A2 => n244, ZN => n92);
   U125 : OR2_X1 port map( A1 => n244, A2 => B(22), ZN => n169);
   U127 : NOR2_X1 port map( A1 => n174, A2 => n99, ZN => n98);
   U129 : NAND2_X1 port map( A1 => B(19), A2 => n247, ZN => n101);
   U130 : NAND2_X1 port map( A1 => n216, A2 => n175, ZN => n173);
   U131 : NOR2_X1 port map( A1 => n247, A2 => B(19), ZN => n102);
   U133 : NAND2_X1 port map( A1 => B(17), A2 => n249, ZN => n107);
   U134 : NAND2_X1 port map( A1 => n175, A2 => n104, ZN => n105);
   U135 : NAND2_X1 port map( A1 => B(18), A2 => n248, ZN => n104);
   U136 : OR2_X1 port map( A1 => n248, A2 => B(18), ZN => n175);
   U138 : NOR2_X1 port map( A1 => n180, A2 => n111, ZN => n110);
   U140 : NAND2_X1 port map( A1 => B(15), A2 => n251, ZN => n113);
   U141 : NAND2_X1 port map( A1 => n220, A2 => n181, ZN => n179);
   U142 : NOR2_X1 port map( A1 => n251, A2 => B(15), ZN => n114);
   U144 : NAND2_X1 port map( A1 => B(13), A2 => n253, ZN => n119);
   U145 : NAND2_X1 port map( A1 => n181, A2 => n116, ZN => n117);
   U146 : NAND2_X1 port map( A1 => B(14), A2 => n252, ZN => n116);
   U147 : OR2_X1 port map( A1 => n252, A2 => B(14), ZN => n181);
   U149 : NOR2_X1 port map( A1 => n186, A2 => n123, ZN => n122);
   U151 : NAND2_X1 port map( A1 => B(11), A2 => n255, ZN => n125);
   U152 : NAND2_X1 port map( A1 => n224, A2 => n187, ZN => n185);
   U153 : NOR2_X1 port map( A1 => n255, A2 => B(11), ZN => n126);
   U155 : NAND2_X1 port map( A1 => B(9), A2 => n257, ZN => n131);
   U156 : NAND2_X1 port map( A1 => n187, A2 => n128, ZN => n129);
   U157 : NAND2_X1 port map( A1 => B(10), A2 => n256, ZN => n128);
   U158 : OR2_X1 port map( A1 => n256, A2 => B(10), ZN => n187);
   U160 : NOR2_X1 port map( A1 => n192, A2 => n135, ZN => n134);
   U162 : NAND2_X1 port map( A1 => B(7), A2 => n259, ZN => n137);
   U163 : NAND2_X1 port map( A1 => n228, A2 => n193, ZN => n191);
   U164 : NOR2_X1 port map( A1 => n259, A2 => B(7), ZN => n138);
   U166 : NAND2_X1 port map( A1 => B(5), A2 => n261, ZN => n143);
   U167 : NAND2_X1 port map( A1 => n193, A2 => n140, ZN => n141);
   U168 : NAND2_X1 port map( A1 => B(6), A2 => n260, ZN => n140);
   U169 : OR2_X1 port map( A1 => n260, A2 => B(6), ZN => n193);
   U171 : NOR2_X1 port map( A1 => n197, A2 => n147, ZN => n146);
   U173 : NAND2_X1 port map( A1 => B(3), A2 => n263, ZN => n149);
   U177 : NAND2_X1 port map( A1 => B(2), A2 => n264, ZN => n153);
   U178 : AOI21_X1 port map( B1 => A(1), B2 => n200, A => n235, ZN => n201);
   U179 : NOR2_X1 port map( A1 => n265, A2 => B(0), ZN => n200);
   U180 : OR2_X1 port map( A1 => n264, A2 => B(2), ZN => n198);
   U181 : NOR2_X1 port map( A1 => n263, A2 => B(3), ZN => n150);
   U182 : NOR2_X1 port map( A1 => n197, A2 => n144, ZN => n194);
   U183 : NOR2_X1 port map( A1 => n261, A2 => B(5), ZN => n144);
   U184 : NOR2_X1 port map( A1 => n262, A2 => B(4), ZN => n197);
   U185 : NOR2_X1 port map( A1 => n192, A2 => n132, ZN => n188);
   U186 : NOR2_X1 port map( A1 => n257, A2 => B(9), ZN => n132);
   U187 : NOR2_X1 port map( A1 => n258, A2 => B(8), ZN => n192);
   U188 : NOR2_X1 port map( A1 => n186, A2 => n120, ZN => n182);
   U189 : NOR2_X1 port map( A1 => n253, A2 => B(13), ZN => n120);
   U190 : NOR2_X1 port map( A1 => n254, A2 => B(12), ZN => n186);
   U191 : NOR2_X1 port map( A1 => n180, A2 => n108, ZN => n176);
   U192 : NOR2_X1 port map( A1 => n249, A2 => B(17), ZN => n108);
   U193 : NOR2_X1 port map( A1 => n250, A2 => B(16), ZN => n180);
   U194 : NOR2_X1 port map( A1 => n174, A2 => n96, ZN => n170);
   U195 : NOR2_X1 port map( A1 => n245, A2 => B(21), ZN => n96);
   U196 : NOR2_X1 port map( A1 => n246, A2 => B(20), ZN => n174);
   U197 : NOR2_X1 port map( A1 => n168, A2 => n84, ZN => n164);
   U198 : NOR2_X1 port map( A1 => n241, A2 => B(25), ZN => n84);
   U199 : NOR2_X1 port map( A1 => n242, A2 => B(24), ZN => n168);
   U200 : NOR2_X1 port map( A1 => n162, A2 => n72, ZN => n158);
   U201 : NOR2_X1 port map( A1 => n237, A2 => B(29), ZN => n72);
   U202 : NOR2_X1 port map( A1 => n238, A2 => B(28), ZN => n162);
   U203 : NOR2_X1 port map( A1 => n204, A2 => A(31), ZN => n66);
   U2 : INV_X1 port map( A => n141, ZN => n229);
   U3 : INV_X1 port map( A => n129, ZN => n225);
   U4 : INV_X1 port map( A => n117, ZN => n221);
   U5 : INV_X1 port map( A => n105, ZN => n217);
   U6 : INV_X1 port map( A => n93, ZN => n213);
   U7 : INV_X1 port map( A => n81, ZN => n209);
   U8 : INV_X1 port map( A => n150, ZN => n232);
   U9 : INV_X1 port map( A => n114, ZN => n220);
   U10 : INV_X1 port map( A => n102, ZN => n216);
   U11 : INV_X1 port map( A => n90, ZN => n212);
   U12 : INV_X1 port map( A => n78, ZN => n208);
   U13 : INV_X1 port map( A => n202, ZN => LE_port);
   U14 : INV_X1 port map( A => n201, ZN => n234);
   U15 : INV_X1 port map( A => A(16), ZN => n250);
   U16 : INV_X1 port map( A => A(15), ZN => n251);
   U17 : INV_X1 port map( A => A(8), ZN => n258);
   U18 : INV_X1 port map( A => A(9), ZN => n257);
   U19 : INV_X1 port map( A => A(5), ZN => n261);
   U20 : INV_X1 port map( A => n138, ZN => n228);
   U21 : INV_X1 port map( A => n126, ZN => n224);
   U22 : INV_X1 port map( A => A(11), ZN => n255);
   U23 : INV_X1 port map( A => A(7), ZN => n259);
   U24 : INV_X1 port map( A => A(6), ZN => n260);
   U25 : INV_X1 port map( A => A(10), ZN => n256);
   U26 : INV_X1 port map( A => A(14), ZN => n252);
   U27 : INV_X1 port map( A => n153, ZN => n233);
   U28 : INV_X1 port map( A => n119, ZN => n223);
   U29 : INV_X1 port map( A => n131, ZN => n227);
   U30 : INV_X1 port map( A => n143, ZN => n231);
   U31 : INV_X1 port map( A => n116, ZN => n222);
   U32 : INV_X1 port map( A => n128, ZN => n226);
   U33 : INV_X1 port map( A => n140, ZN => n230);
   U34 : INV_X1 port map( A => A(28), ZN => n238);
   U35 : INV_X1 port map( A => A(17), ZN => n249);
   U36 : INV_X1 port map( A => A(21), ZN => n245);
   U37 : INV_X1 port map( A => A(25), ZN => n241);
   U38 : INV_X1 port map( A => A(20), ZN => n246);
   U39 : INV_X1 port map( A => A(27), ZN => n239);
   U40 : INV_X1 port map( A => A(19), ZN => n247);
   U41 : INV_X1 port map( A => A(26), ZN => n240);
   U42 : INV_X1 port map( A => n83, ZN => n211);
   U43 : INV_X1 port map( A => n80, ZN => n210);
   U44 : INV_X1 port map( A => n95, ZN => n215);
   U45 : INV_X1 port map( A => n107, ZN => n219);
   U46 : INV_X1 port map( A => n104, ZN => n218);
   U47 : INV_X1 port map( A => n92, ZN => n214);
   U48 : INV_X1 port map( A => n71, ZN => n207);
   U49 : INV_X1 port map( A => n67, ZN => n205);
   U50 : INV_X1 port map( A => A(30), ZN => n236);
   U51 : INV_X1 port map( A => A(13), ZN => n253);
   U52 : INV_X1 port map( A => A(12), ZN => n254);
   U53 : INV_X1 port map( A => A(4), ZN => n262);
   U54 : INV_X1 port map( A => B(1), ZN => n235);
   U55 : INV_X1 port map( A => A(3), ZN => n263);
   U56 : INV_X1 port map( A => A(2), ZN => n264);
   U57 : INV_X1 port map( A => A(24), ZN => n242);
   U58 : INV_X1 port map( A => A(29), ZN => n237);
   U59 : INV_X1 port map( A => A(23), ZN => n243);
   U60 : INV_X1 port map( A => A(18), ZN => n248);
   U61 : INV_X1 port map( A => A(22), ZN => n244);
   U62 : INV_X1 port map( A => B(30), ZN => n206);
   U63 : INV_X1 port map( A => B(31), ZN => n204);
   U64 : INV_X1 port map( A => A(0), ZN => n265);
   U1 : OAI211_X1 port map( C1 => n190, C2 => n191, A => n137, B => n134, ZN =>
                           n189);
   U104 : AOI211_X1 port map( C1 => n194, C2 => n195, A => n141, B => n231, ZN 
                           => n190);
   U106 : OAI211_X1 port map( C1 => n178, C2 => n179, A => n113, B => n110, ZN 
                           => n177);
   U110 : AOI211_X1 port map( C1 => n182, C2 => n183, A => n117, B => n223, ZN 
                           => n178);
   U115 : OAI211_X1 port map( C1 => n166, C2 => n167, A => n89, B => n86, ZN =>
                           n165);
   U117 : AOI211_X1 port map( C1 => n170, C2 => n171, A => n93, B => n215, ZN 
                           => n166);
   U121 : NAND3_X1 port map( A1 => n196, A2 => n149, A3 => n146, ZN => n195);
   U126 : NAND3_X1 port map( A1 => n232, A2 => n198, A3 => n199, ZN => n196);
   U128 : OAI211_X1 port map( C1 => A(1), C2 => n200, A => n234, B => n152, ZN 
                           => n199);
   U132 : AND2_X1 port map( A1 => B(4), A2 => n262, ZN => n147);
   U137 : AND2_X1 port map( A1 => n198, A2 => n153, ZN => n152);
   U139 : AND2_X1 port map( A1 => B(8), A2 => n258, ZN => n135);
   U143 : OAI211_X1 port map( C1 => n184, C2 => n185, A => n125, B => n122, ZN 
                           => n183);
   U148 : AOI211_X1 port map( C1 => n188, C2 => n189, A => n129, B => n227, ZN 
                           => n184);
   U150 : AND2_X1 port map( A1 => B(12), A2 => n254, ZN => n123);
   U154 : AND2_X1 port map( A1 => B(16), A2 => n250, ZN => n111);
   U159 : OAI211_X1 port map( C1 => n172, C2 => n173, A => n101, B => n98, ZN 
                           => n171);
   U161 : AOI211_X1 port map( C1 => n176, C2 => n177, A => n105, B => n219, ZN 
                           => n172);
   U165 : AND2_X1 port map( A1 => B(20), A2 => n246, ZN => n99);
   U170 : AND2_X1 port map( A1 => B(24), A2 => n242, ZN => n87);
   U172 : OAI211_X1 port map( C1 => n160, C2 => n161, A => n77, B => n74, ZN =>
                           n159);
   U174 : AOI211_X1 port map( C1 => n164, C2 => n165, A => n81, B => n211, ZN 
                           => n160);
   U175 : AND2_X1 port map( A1 => B(28), A2 => n238, ZN => n75);
   U176 : AND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => EQ);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end ALU_N32_DW01_cmp6_0;

architecture SYN_rpl of ALU_N32_DW01_cmp6_0 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n202, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78
      , n79, n81, n82, n84, n85, n86, n87, n88, n89, n91, n92, n94, n95, n96, 
      n97, n98, n99, n101, n102, n104, n105, n106, n107, n108, n109, n111, n112
      , n114, n115, n116, n117, n118, n119, n121, n122, n124, n125, n126, n127,
      n128, n129, n131, n132, n134, n135, n136, n137, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n93, n90, n83
      , n80, n73, n200, n138, n133, n130, n123, n120, n113, n110, n103, n100, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266 : std_logic;

begin
   
   U65 : AOI21_X1 port map( B1 => n65, B2 => n205, A => n66, ZN => LE);
   U66 : AOI22_X1 port map( A1 => A(30), A2 => n206, B1 => n68, B2 => n69, ZN 
                           => n67);
   U67 : AOI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n68);
   U69 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n74);
   U72 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n84);
   U75 : NAND2_X1 port map( A1 => n97, A2 => n98, ZN => n94);
   U78 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => n104);
   U81 : NAND2_X1 port map( A1 => n117, A2 => n118, ZN => n114);
   U84 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => n124);
   U89 : OAI21_X1 port map( B1 => n266, B2 => n141, A => B(1), ZN => n139);
   U90 : NAND2_X1 port map( A1 => A(0), A2 => n264, ZN => n141);
   U91 : NOR2_X1 port map( A1 => n142, A2 => n143, ZN => n129);
   U92 : NOR2_X1 port map( A1 => n144, A2 => n145, ZN => n119);
   U93 : NOR2_X1 port map( A1 => n146, A2 => n147, ZN => n109);
   U94 : NOR2_X1 port map( A1 => n148, A2 => n149, ZN => n99);
   U95 : NOR2_X1 port map( A1 => n150, A2 => n151, ZN => n89);
   U96 : NOR2_X1 port map( A1 => n152, A2 => n153, ZN => n79);
   U97 : NOR2_X1 port map( A1 => n154, A2 => n155, ZN => n70);
   U98 : OAI21_X1 port map( B1 => n66, B2 => n156, A => n65, ZN => n202);
   U99 : NAND2_X1 port map( A1 => A(31), A2 => n204, ZN => n65);
   U100 : AOI22_X1 port map( A1 => B(30), A2 => n265, B1 => n157, B2 => n69, ZN
                           => n156);
   U101 : XOR2_X1 port map( A => n265, B => B(30), Z => n69);
   U102 : AOI21_X1 port map( B1 => n158, B2 => n207, A => n155, ZN => n157);
   U104 : NOR2_X1 port map( A1 => n208, A2 => A(29), ZN => n72);
   U105 : AOI21_X1 port map( B1 => n159, B2 => n76, A => n160, ZN => n158);
   U106 : NOR2_X1 port map( A1 => n160, A2 => n154, ZN => n76);
   U108 : NOR2_X1 port map( A1 => n209, A2 => A(28), ZN => n160);
   U109 : AOI21_X1 port map( B1 => n161, B2 => n75, A => n210, ZN => n159);
   U110 : NAND2_X1 port map( A1 => A(27), A2 => n211, ZN => n77);
   U111 : OR2_X1 port map( A1 => n211, A2 => A(27), ZN => n75);
   U112 : AOI21_X1 port map( B1 => n162, B2 => n212, A => n163, ZN => n161);
   U113 : NAND2_X1 port map( A1 => n213, A2 => n78, ZN => n81);
   U114 : NAND2_X1 port map( A1 => A(26), A2 => n214, ZN => n78);
   U115 : NOR2_X1 port map( A1 => n214, A2 => A(26), ZN => n163);
   U116 : AOI21_X1 port map( B1 => n164, B2 => n215, A => n153, ZN => n162);
   U118 : NOR2_X1 port map( A1 => n216, A2 => A(25), ZN => n82);
   U119 : AOI21_X1 port map( B1 => n165, B2 => n86, A => n166, ZN => n164);
   U120 : NOR2_X1 port map( A1 => n166, A2 => n152, ZN => n86);
   U122 : NOR2_X1 port map( A1 => n217, A2 => A(24), ZN => n166);
   U123 : AOI21_X1 port map( B1 => n167, B2 => n85, A => n218, ZN => n165);
   U124 : NAND2_X1 port map( A1 => A(23), A2 => n219, ZN => n87);
   U125 : OR2_X1 port map( A1 => n219, A2 => A(23), ZN => n85);
   U126 : AOI21_X1 port map( B1 => n168, B2 => n220, A => n169, ZN => n167);
   U127 : NAND2_X1 port map( A1 => n221, A2 => n88, ZN => n91);
   U128 : NAND2_X1 port map( A1 => A(22), A2 => n222, ZN => n88);
   U129 : NOR2_X1 port map( A1 => n222, A2 => A(22), ZN => n169);
   U130 : AOI21_X1 port map( B1 => n170, B2 => n223, A => n151, ZN => n168);
   U132 : NOR2_X1 port map( A1 => n224, A2 => A(21), ZN => n92);
   U133 : AOI21_X1 port map( B1 => n171, B2 => n96, A => n172, ZN => n170);
   U134 : NOR2_X1 port map( A1 => n172, A2 => n150, ZN => n96);
   U136 : NOR2_X1 port map( A1 => n225, A2 => A(20), ZN => n172);
   U137 : AOI21_X1 port map( B1 => n173, B2 => n95, A => n226, ZN => n171);
   U138 : NAND2_X1 port map( A1 => A(19), A2 => n227, ZN => n97);
   U139 : OR2_X1 port map( A1 => n227, A2 => A(19), ZN => n95);
   U140 : AOI21_X1 port map( B1 => n174, B2 => n228, A => n175, ZN => n173);
   U141 : NAND2_X1 port map( A1 => n229, A2 => n98, ZN => n101);
   U142 : NAND2_X1 port map( A1 => A(18), A2 => n230, ZN => n98);
   U143 : NOR2_X1 port map( A1 => n230, A2 => A(18), ZN => n175);
   U144 : AOI21_X1 port map( B1 => n176, B2 => n231, A => n149, ZN => n174);
   U146 : NOR2_X1 port map( A1 => n232, A2 => A(17), ZN => n102);
   U147 : AOI21_X1 port map( B1 => n177, B2 => n106, A => n178, ZN => n176);
   U148 : NOR2_X1 port map( A1 => n178, A2 => n148, ZN => n106);
   U150 : NOR2_X1 port map( A1 => n233, A2 => A(16), ZN => n178);
   U151 : AOI21_X1 port map( B1 => n179, B2 => n105, A => n234, ZN => n177);
   U152 : NAND2_X1 port map( A1 => A(15), A2 => n235, ZN => n107);
   U153 : OR2_X1 port map( A1 => n235, A2 => A(15), ZN => n105);
   U154 : AOI21_X1 port map( B1 => n180, B2 => n236, A => n181, ZN => n179);
   U155 : NAND2_X1 port map( A1 => n237, A2 => n108, ZN => n111);
   U156 : NAND2_X1 port map( A1 => A(14), A2 => n238, ZN => n108);
   U157 : NOR2_X1 port map( A1 => n238, A2 => A(14), ZN => n181);
   U158 : AOI21_X1 port map( B1 => n182, B2 => n239, A => n147, ZN => n180);
   U160 : NOR2_X1 port map( A1 => n240, A2 => A(13), ZN => n112);
   U161 : AOI21_X1 port map( B1 => n183, B2 => n116, A => n184, ZN => n182);
   U162 : NOR2_X1 port map( A1 => n184, A2 => n146, ZN => n116);
   U164 : NOR2_X1 port map( A1 => n241, A2 => A(12), ZN => n184);
   U165 : AOI21_X1 port map( B1 => n185, B2 => n115, A => n242, ZN => n183);
   U166 : NAND2_X1 port map( A1 => A(11), A2 => n243, ZN => n117);
   U167 : OR2_X1 port map( A1 => n243, A2 => A(11), ZN => n115);
   U168 : AOI21_X1 port map( B1 => n186, B2 => n244, A => n187, ZN => n185);
   U169 : NAND2_X1 port map( A1 => n245, A2 => n118, ZN => n121);
   U170 : NAND2_X1 port map( A1 => A(10), A2 => n246, ZN => n118);
   U171 : NOR2_X1 port map( A1 => n246, A2 => A(10), ZN => n187);
   U172 : AOI21_X1 port map( B1 => n188, B2 => n247, A => n145, ZN => n186);
   U174 : NOR2_X1 port map( A1 => n248, A2 => A(9), ZN => n122);
   U175 : AOI21_X1 port map( B1 => n189, B2 => n126, A => n190, ZN => n188);
   U176 : NOR2_X1 port map( A1 => n190, A2 => n144, ZN => n126);
   U178 : NOR2_X1 port map( A1 => n249, A2 => A(8), ZN => n190);
   U179 : AOI21_X1 port map( B1 => n191, B2 => n125, A => n250, ZN => n189);
   U180 : NAND2_X1 port map( A1 => A(7), A2 => n251, ZN => n127);
   U181 : OR2_X1 port map( A1 => n251, A2 => A(7), ZN => n125);
   U182 : AOI21_X1 port map( B1 => n192, B2 => n252, A => n193, ZN => n191);
   U183 : NAND2_X1 port map( A1 => n253, A2 => n128, ZN => n131);
   U184 : NAND2_X1 port map( A1 => A(6), A2 => n254, ZN => n128);
   U185 : NOR2_X1 port map( A1 => n254, A2 => A(6), ZN => n193);
   U186 : AOI21_X1 port map( B1 => n194, B2 => n255, A => n143, ZN => n192);
   U188 : NOR2_X1 port map( A1 => n256, A2 => A(5), ZN => n132);
   U189 : AOI21_X1 port map( B1 => n195, B2 => n135, A => n196, ZN => n194);
   U190 : NOR2_X1 port map( A1 => n196, A2 => n142, ZN => n135);
   U192 : NOR2_X1 port map( A1 => n257, A2 => A(4), ZN => n196);
   U193 : AOI21_X1 port map( B1 => n197, B2 => n134, A => n258, ZN => n195);
   U194 : NAND2_X1 port map( A1 => A(3), A2 => n259, ZN => n136);
   U195 : OR2_X1 port map( A1 => n259, A2 => A(3), ZN => n134);
   U196 : AOI21_X1 port map( B1 => n262, B2 => n140, A => n198, ZN => n197);
   U197 : NOR2_X1 port map( A1 => n198, A2 => n260, ZN => n140);
   U198 : NAND2_X1 port map( A1 => A(2), A2 => n261, ZN => n137);
   U199 : NOR2_X1 port map( A1 => n261, A2 => A(2), ZN => n198);
   U202 : NOR2_X1 port map( A1 => n264, A2 => A(0), ZN => n201);
   U203 : NOR2_X1 port map( A1 => n204, A2 => A(31), ZN => n66);
   U1 : INV_X1 port map( A => n121, ZN => n244);
   U2 : INV_X1 port map( A => n81, ZN => n212);
   U3 : INV_X1 port map( A => n131, ZN => n252);
   U4 : INV_X1 port map( A => n132, ZN => n255);
   U5 : INV_X1 port map( A => n77, ZN => n210);
   U6 : INV_X1 port map( A => n122, ZN => n247);
   U7 : INV_X1 port map( A => n102, ZN => n231);
   U8 : INV_X1 port map( A => n193, ZN => n253);
   U9 : INV_X1 port map( A => n181, ZN => n237);
   U10 : INV_X1 port map( A => n187, ZN => n245);
   U11 : INV_X1 port map( A => n127, ZN => n250);
   U12 : INV_X1 port map( A => n163, ZN => n213);
   U13 : INV_X1 port map( A => n101, ZN => n228);
   U14 : INV_X1 port map( A => n107, ZN => n234);
   U15 : INV_X1 port map( A => n137, ZN => n260);
   U16 : INV_X1 port map( A => n136, ZN => n258);
   U17 : INV_X1 port map( A => n117, ZN => n242);
   U18 : INV_X1 port map( A => n91, ZN => n220);
   U19 : INV_X1 port map( A => n92, ZN => n223);
   U20 : INV_X1 port map( A => n111, ZN => n236);
   U21 : INV_X1 port map( A => n112, ZN => n239);
   U22 : INV_X1 port map( A => n97, ZN => n226);
   U23 : INV_X1 port map( A => n82, ZN => n215);
   U24 : INV_X1 port map( A => A(1), ZN => n266);
   U25 : INV_X1 port map( A => B(4), ZN => n257);
   U26 : INV_X1 port map( A => n67, ZN => n205);
   U27 : INV_X1 port map( A => n175, ZN => n229);
   U28 : INV_X1 port map( A => n169, ZN => n221);
   U29 : INV_X1 port map( A => A(30), ZN => n265);
   U30 : INV_X1 port map( A => n72, ZN => n207);
   U31 : INV_X1 port map( A => n87, ZN => n218);
   U32 : INV_X1 port map( A => n141, ZN => n263);
   U33 : INV_X1 port map( A => B(0), ZN => n264);
   U34 : INV_X1 port map( A => B(3), ZN => n259);
   U35 : INV_X1 port map( A => B(2), ZN => n261);
   U36 : INV_X1 port map( A => B(9), ZN => n248);
   U37 : INV_X1 port map( A => B(12), ZN => n241);
   U38 : INV_X1 port map( A => B(14), ZN => n238);
   U39 : INV_X1 port map( A => B(8), ZN => n249);
   U40 : INV_X1 port map( A => B(5), ZN => n256);
   U41 : INV_X1 port map( A => B(10), ZN => n246);
   U42 : INV_X1 port map( A => B(6), ZN => n254);
   U43 : INV_X1 port map( A => B(11), ZN => n243);
   U44 : INV_X1 port map( A => n202, ZN => GE);
   U45 : INV_X1 port map( A => B(7), ZN => n251);
   U46 : INV_X1 port map( A => n199, ZN => n262);
   U47 : INV_X1 port map( A => B(13), ZN => n240);
   U48 : INV_X1 port map( A => B(28), ZN => n209);
   U49 : INV_X1 port map( A => B(25), ZN => n216);
   U50 : INV_X1 port map( A => B(26), ZN => n214);
   U51 : INV_X1 port map( A => B(31), ZN => n204);
   U52 : INV_X1 port map( A => B(21), ZN => n224);
   U53 : INV_X1 port map( A => B(20), ZN => n225);
   U54 : INV_X1 port map( A => B(17), ZN => n232);
   U55 : INV_X1 port map( A => B(16), ZN => n233);
   U56 : INV_X1 port map( A => B(18), ZN => n230);
   U57 : INV_X1 port map( A => B(29), ZN => n208);
   U58 : INV_X1 port map( A => B(24), ZN => n217);
   U59 : INV_X1 port map( A => B(22), ZN => n222);
   U60 : INV_X1 port map( A => B(27), ZN => n211);
   U61 : INV_X1 port map( A => B(19), ZN => n227);
   U62 : INV_X1 port map( A => B(23), ZN => n219);
   U63 : INV_X1 port map( A => B(30), ZN => n206);
   U64 : INV_X1 port map( A => B(15), ZN => n235);
   U68 : AND2_X1 port map( A1 => A(4), A2 => n257, ZN => n142);
   U70 : AND2_X1 port map( A1 => A(5), A2 => n256, ZN => n143);
   U71 : OAI211_X1 port map( C1 => A(1), C2 => n263, A => n139, B => n140, ZN 
                           => n138);
   U73 : AND2_X1 port map( A1 => A(13), A2 => n240, ZN => n147);
   U74 : AND2_X1 port map( A1 => A(12), A2 => n241, ZN => n146);
   U76 : AOI211_X1 port map( C1 => n119, C2 => n120, A => n121, B => n122, ZN 
                           => n113);
   U77 : OAI211_X1 port map( C1 => n123, C2 => n124, A => n125, B => n126, ZN 
                           => n120);
   U79 : AND2_X1 port map( A1 => A(20), A2 => n225, ZN => n150);
   U80 : AOI211_X1 port map( C1 => n99, C2 => n100, A => n101, B => n102, ZN =>
                           n93);
   U82 : OAI211_X1 port map( C1 => n103, C2 => n104, A => n105, B => n106, ZN 
                           => n100);
   U83 : AOI211_X1 port map( C1 => n79, C2 => n80, A => n81, B => n82, ZN => 
                           n73);
   U85 : OAI211_X1 port map( C1 => n83, C2 => n84, A => n85, B => n86, ZN => 
                           n80);
   U86 : OAI22_X1 port map( A1 => n200, A2 => B(1), B1 => n266, B2 => n201, ZN 
                           => n199);
   U87 : AND2_X1 port map( A1 => n201, A2 => n266, ZN => n200);
   U88 : AND2_X1 port map( A1 => A(9), A2 => n248, ZN => n145);
   U103 : AND2_X1 port map( A1 => A(8), A2 => n249, ZN => n144);
   U107 : AOI211_X1 port map( C1 => n129, C2 => n130, A => n131, B => n132, ZN 
                           => n123);
   U117 : NAND3_X1 port map( A1 => n133, A2 => n134, A3 => n135, ZN => n130);
   U121 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n138, ZN => n133);
   U131 : AND2_X1 port map( A1 => A(17), A2 => n232, ZN => n149);
   U135 : AND2_X1 port map( A1 => A(16), A2 => n233, ZN => n148);
   U145 : AOI211_X1 port map( C1 => n109, C2 => n110, A => n111, B => n112, ZN 
                           => n103);
   U149 : OAI211_X1 port map( C1 => n113, C2 => n114, A => n115, B => n116, ZN 
                           => n110);
   U159 : AND2_X1 port map( A1 => A(21), A2 => n224, ZN => n151);
   U163 : AND2_X1 port map( A1 => A(24), A2 => n217, ZN => n152);
   U173 : AND2_X1 port map( A1 => A(25), A2 => n216, ZN => n153);
   U177 : AOI211_X1 port map( C1 => n89, C2 => n90, A => n91, B => n92, ZN => 
                           n83);
   U187 : OAI211_X1 port map( C1 => n93, C2 => n94, A => n95, B => n96, ZN => 
                           n90);
   U191 : AND2_X1 port map( A1 => A(28), A2 => n209, ZN => n154);
   U200 : AND2_X1 port map( A1 => A(29), A2 => n208, ZN => n155);
   U201 : OAI211_X1 port map( C1 => n73, C2 => n74, A => n75, B => n76, ZN => 
                           n71);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity pc_add_N32_OP24_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end pc_add_N32_OP24_DW01_add_0;

architecture SYN_rpl of pc_add_N32_OP24_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, SUM_7_port, 
      SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port, 
      SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, SUM_31_port, n30, n31, n32, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      , n49, n50, n51, n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U2 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U3 : XOR2_X1 port map( A => A(4), B => n30, Z => SUM_4_port);
   U4 : XOR2_X1 port map( A => A(5), B => n31, Z => SUM_5_port);
   U5 : XOR2_X1 port map( A => A(6), B => n32, Z => SUM_6_port);
   U6 : XOR2_X1 port map( A => A(7), B => n33, Z => SUM_7_port);
   U7 : XOR2_X1 port map( A => A(8), B => n34, Z => SUM_8_port);
   U8 : XOR2_X1 port map( A => A(9), B => n35, Z => SUM_9_port);
   U9 : XOR2_X1 port map( A => A(10), B => n36, Z => SUM_10_port);
   U10 : XOR2_X1 port map( A => A(11), B => n37, Z => SUM_11_port);
   U11 : XOR2_X1 port map( A => A(12), B => n38, Z => SUM_12_port);
   U12 : XOR2_X1 port map( A => A(13), B => n39, Z => SUM_13_port);
   U13 : XOR2_X1 port map( A => A(14), B => n40, Z => SUM_14_port);
   U14 : XOR2_X1 port map( A => A(15), B => n41, Z => SUM_15_port);
   U15 : XOR2_X1 port map( A => A(16), B => n42, Z => SUM_16_port);
   U16 : XOR2_X1 port map( A => A(17), B => n43, Z => SUM_17_port);
   U17 : XOR2_X1 port map( A => A(18), B => n44, Z => SUM_18_port);
   U18 : XOR2_X1 port map( A => A(19), B => n45, Z => SUM_19_port);
   U19 : XOR2_X1 port map( A => A(20), B => n46, Z => SUM_20_port);
   U20 : XOR2_X1 port map( A => A(21), B => n47, Z => SUM_21_port);
   U21 : XOR2_X1 port map( A => A(22), B => n48, Z => SUM_22_port);
   U22 : XOR2_X1 port map( A => A(23), B => n49, Z => SUM_23_port);
   U23 : XOR2_X1 port map( A => A(24), B => n50, Z => SUM_24_port);
   U24 : XOR2_X1 port map( A => A(25), B => n51, Z => SUM_25_port);
   U25 : XOR2_X1 port map( A => A(26), B => n52, Z => SUM_26_port);
   U26 : XOR2_X1 port map( A => A(27), B => n53, Z => SUM_27_port);
   U27 : XOR2_X1 port map( A => A(28), B => n54, Z => SUM_28_port);
   U28 : XOR2_X1 port map( A => A(29), B => n55, Z => SUM_29_port);
   U29 : XOR2_X1 port map( A => A(30), B => n56, Z => SUM_30_port);
   U30 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U58 : NAND2_X1 port map( A1 => A(30), A2 => n56, ZN => n57);
   U1 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U31 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n30);
   U32 : AND2_X1 port map( A1 => A(4), A2 => n30, ZN => n31);
   U33 : AND2_X1 port map( A1 => A(5), A2 => n31, ZN => n32);
   U34 : AND2_X1 port map( A1 => A(6), A2 => n32, ZN => n33);
   U35 : AND2_X1 port map( A1 => A(7), A2 => n33, ZN => n34);
   U36 : AND2_X1 port map( A1 => A(8), A2 => n34, ZN => n35);
   U37 : AND2_X1 port map( A1 => A(9), A2 => n35, ZN => n36);
   U38 : AND2_X1 port map( A1 => A(10), A2 => n36, ZN => n37);
   U39 : AND2_X1 port map( A1 => A(11), A2 => n37, ZN => n38);
   U40 : AND2_X1 port map( A1 => A(12), A2 => n38, ZN => n39);
   U41 : AND2_X1 port map( A1 => A(13), A2 => n39, ZN => n40);
   U42 : AND2_X1 port map( A1 => A(14), A2 => n40, ZN => n41);
   U43 : AND2_X1 port map( A1 => A(15), A2 => n41, ZN => n42);
   U44 : AND2_X1 port map( A1 => A(16), A2 => n42, ZN => n43);
   U45 : AND2_X1 port map( A1 => A(17), A2 => n43, ZN => n44);
   U46 : AND2_X1 port map( A1 => A(18), A2 => n44, ZN => n45);
   U47 : AND2_X1 port map( A1 => A(19), A2 => n45, ZN => n46);
   U48 : AND2_X1 port map( A1 => A(20), A2 => n46, ZN => n47);
   U49 : AND2_X1 port map( A1 => A(21), A2 => n47, ZN => n48);
   U50 : AND2_X1 port map( A1 => A(22), A2 => n48, ZN => n49);
   U51 : AND2_X1 port map( A1 => A(23), A2 => n49, ZN => n50);
   U52 : AND2_X1 port map( A1 => A(24), A2 => n50, ZN => n51);
   U53 : AND2_X1 port map( A1 => A(25), A2 => n51, ZN => n52);
   U54 : AND2_X1 port map( A1 => A(26), A2 => n52, ZN => n53);
   U55 : AND2_X1 port map( A1 => A(27), A2 => n53, ZN => n54);
   U56 : AND2_X1 port map( A1 => A(28), A2 => n54, ZN => n55);
   U57 : AND2_X1 port map( A1 => A(29), A2 => n55, ZN => n56);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_mux41_N32 is

   port( sel : in std_logic_vector (1 downto 0);  w, x, y, z : in 
         std_logic_vector (31 downto 0);  m : out std_logic_vector (31 downto 
         0));

end gen_mux41_N32;

architecture SYN_dflow of gen_mux41_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n74, n77, n80, n83, n84, 
      n85 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => m(9));
   U4 : AOI22_X1 port map( A1 => w(9), A2 => n83, B1 => x(9), B2 => n80, ZN => 
                           n4);
   U5 : AOI22_X1 port map( A1 => y(9), A2 => n77, B1 => z(9), B2 => n74, ZN => 
                           n3);
   U6 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => m(8));
   U7 : AOI22_X1 port map( A1 => w(8), A2 => n83, B1 => x(8), B2 => n80, ZN => 
                           n10);
   U8 : AOI22_X1 port map( A1 => y(8), A2 => n77, B1 => z(8), B2 => n74, ZN => 
                           n9);
   U9 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => m(7));
   U10 : AOI22_X1 port map( A1 => w(7), A2 => n83, B1 => x(7), B2 => n80, ZN =>
                           n12);
   U11 : AOI22_X1 port map( A1 => y(7), A2 => n77, B1 => z(7), B2 => n74, ZN =>
                           n11);
   U12 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => m(6));
   U13 : AOI22_X1 port map( A1 => w(6), A2 => n83, B1 => x(6), B2 => n80, ZN =>
                           n14);
   U14 : AOI22_X1 port map( A1 => y(6), A2 => n77, B1 => z(6), B2 => n74, ZN =>
                           n13);
   U15 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => m(5));
   U16 : AOI22_X1 port map( A1 => w(5), A2 => n83, B1 => x(5), B2 => n80, ZN =>
                           n16);
   U17 : AOI22_X1 port map( A1 => y(5), A2 => n77, B1 => z(5), B2 => n74, ZN =>
                           n15);
   U18 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => m(4));
   U19 : AOI22_X1 port map( A1 => w(4), A2 => n83, B1 => x(4), B2 => n80, ZN =>
                           n18);
   U20 : AOI22_X1 port map( A1 => y(4), A2 => n77, B1 => z(4), B2 => n74, ZN =>
                           n17);
   U21 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => m(3));
   U22 : AOI22_X1 port map( A1 => w(3), A2 => n83, B1 => x(3), B2 => n80, ZN =>
                           n20);
   U23 : AOI22_X1 port map( A1 => y(3), A2 => n77, B1 => z(3), B2 => n74, ZN =>
                           n19);
   U24 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => m(31));
   U25 : AOI22_X1 port map( A1 => w(31), A2 => n83, B1 => x(31), B2 => n80, ZN 
                           => n22);
   U26 : AOI22_X1 port map( A1 => y(31), A2 => n77, B1 => z(31), B2 => n74, ZN 
                           => n21);
   U27 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => m(30));
   U28 : AOI22_X1 port map( A1 => w(30), A2 => n83, B1 => x(30), B2 => n6, ZN 
                           => n24);
   U29 : AOI22_X1 port map( A1 => y(30), A2 => n77, B1 => z(30), B2 => n8, ZN 
                           => n23);
   U30 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => m(2));
   U31 : AOI22_X1 port map( A1 => w(2), A2 => n5, B1 => x(2), B2 => n80, ZN => 
                           n26);
   U32 : AOI22_X1 port map( A1 => y(2), A2 => n7, B1 => z(2), B2 => n74, ZN => 
                           n25);
   U33 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => m(29));
   U34 : AOI22_X1 port map( A1 => w(29), A2 => n83, B1 => x(29), B2 => n80, ZN 
                           => n28);
   U35 : AOI22_X1 port map( A1 => y(29), A2 => n77, B1 => z(29), B2 => n8, ZN 
                           => n27);
   U36 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => m(28));
   U37 : AOI22_X1 port map( A1 => w(28), A2 => n83, B1 => x(28), B2 => n6, ZN 
                           => n30);
   U38 : AOI22_X1 port map( A1 => y(28), A2 => n77, B1 => z(28), B2 => n8, ZN 
                           => n29);
   U39 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => m(27));
   U40 : AOI22_X1 port map( A1 => w(27), A2 => n83, B1 => x(27), B2 => n80, ZN 
                           => n32);
   U41 : AOI22_X1 port map( A1 => y(27), A2 => n7, B1 => z(27), B2 => n74, ZN 
                           => n31);
   U42 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => m(26));
   U43 : AOI22_X1 port map( A1 => w(26), A2 => n83, B1 => x(26), B2 => n80, ZN 
                           => n34);
   U44 : AOI22_X1 port map( A1 => y(26), A2 => n7, B1 => z(26), B2 => n74, ZN 
                           => n33);
   U45 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => m(25));
   U46 : AOI22_X1 port map( A1 => w(25), A2 => n5, B1 => x(25), B2 => n80, ZN 
                           => n36);
   U47 : AOI22_X1 port map( A1 => y(25), A2 => n7, B1 => z(25), B2 => n74, ZN 
                           => n35);
   U48 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => m(24));
   U49 : AOI22_X1 port map( A1 => w(24), A2 => n83, B1 => x(24), B2 => n80, ZN 
                           => n38);
   U50 : AOI22_X1 port map( A1 => y(24), A2 => n77, B1 => z(24), B2 => n74, ZN 
                           => n37);
   U51 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => m(23));
   U52 : AOI22_X1 port map( A1 => w(23), A2 => n83, B1 => x(23), B2 => n80, ZN 
                           => n40);
   U53 : AOI22_X1 port map( A1 => y(23), A2 => n77, B1 => z(23), B2 => n8, ZN 
                           => n39);
   U54 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => m(22));
   U55 : AOI22_X1 port map( A1 => w(22), A2 => n83, B1 => x(22), B2 => n80, ZN 
                           => n42);
   U56 : AOI22_X1 port map( A1 => y(22), A2 => n77, B1 => z(22), B2 => n74, ZN 
                           => n41);
   U57 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => m(21));
   U58 : AOI22_X1 port map( A1 => w(21), A2 => n5, B1 => x(21), B2 => n80, ZN 
                           => n44);
   U59 : AOI22_X1 port map( A1 => y(21), A2 => n7, B1 => z(21), B2 => n74, ZN 
                           => n43);
   U60 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => m(20));
   U61 : AOI22_X1 port map( A1 => w(20), A2 => n83, B1 => x(20), B2 => n6, ZN 
                           => n46);
   U62 : AOI22_X1 port map( A1 => y(20), A2 => n77, B1 => z(20), B2 => n74, ZN 
                           => n45);
   U63 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => m(1));
   U64 : AOI22_X1 port map( A1 => w(1), A2 => n5, B1 => x(1), B2 => n6, ZN => 
                           n48);
   U65 : AOI22_X1 port map( A1 => y(1), A2 => n7, B1 => z(1), B2 => n8, ZN => 
                           n47);
   U66 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => m(19));
   U67 : AOI22_X1 port map( A1 => w(19), A2 => n5, B1 => x(19), B2 => n6, ZN =>
                           n50);
   U68 : AOI22_X1 port map( A1 => y(19), A2 => n77, B1 => z(19), B2 => n8, ZN 
                           => n49);
   U69 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => m(18));
   U70 : AOI22_X1 port map( A1 => w(18), A2 => n5, B1 => x(18), B2 => n6, ZN =>
                           n52);
   U71 : AOI22_X1 port map( A1 => y(18), A2 => n7, B1 => z(18), B2 => n8, ZN =>
                           n51);
   U72 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => m(17));
   U73 : AOI22_X1 port map( A1 => w(17), A2 => n83, B1 => x(17), B2 => n80, ZN 
                           => n54);
   U74 : AOI22_X1 port map( A1 => y(17), A2 => n77, B1 => z(17), B2 => n74, ZN 
                           => n53);
   U75 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => m(16));
   U76 : AOI22_X1 port map( A1 => w(16), A2 => n83, B1 => x(16), B2 => n80, ZN 
                           => n56);
   U77 : AOI22_X1 port map( A1 => y(16), A2 => n77, B1 => z(16), B2 => n74, ZN 
                           => n55);
   U78 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => m(15));
   U79 : AOI22_X1 port map( A1 => w(15), A2 => n83, B1 => x(15), B2 => n80, ZN 
                           => n58);
   U80 : AOI22_X1 port map( A1 => y(15), A2 => n77, B1 => z(15), B2 => n74, ZN 
                           => n57);
   U81 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => m(14));
   U82 : AOI22_X1 port map( A1 => w(14), A2 => n83, B1 => x(14), B2 => n80, ZN 
                           => n60);
   U83 : AOI22_X1 port map( A1 => y(14), A2 => n77, B1 => z(14), B2 => n74, ZN 
                           => n59);
   U84 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => m(13));
   U85 : AOI22_X1 port map( A1 => w(13), A2 => n5, B1 => x(13), B2 => n6, ZN =>
                           n62);
   U86 : AOI22_X1 port map( A1 => y(13), A2 => n7, B1 => z(13), B2 => n8, ZN =>
                           n61);
   U87 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => m(12));
   U88 : AOI22_X1 port map( A1 => w(12), A2 => n5, B1 => x(12), B2 => n6, ZN =>
                           n64);
   U89 : AOI22_X1 port map( A1 => y(12), A2 => n7, B1 => z(12), B2 => n8, ZN =>
                           n63);
   U90 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => m(11));
   U91 : AOI22_X1 port map( A1 => w(11), A2 => n5, B1 => x(11), B2 => n6, ZN =>
                           n66);
   U92 : AOI22_X1 port map( A1 => y(11), A2 => n7, B1 => z(11), B2 => n8, ZN =>
                           n65);
   U93 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => m(10));
   U94 : AOI22_X1 port map( A1 => w(10), A2 => n5, B1 => x(10), B2 => n6, ZN =>
                           n68);
   U95 : AOI22_X1 port map( A1 => y(10), A2 => n7, B1 => z(10), B2 => n8, ZN =>
                           n67);
   U96 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => m(0));
   U97 : AOI22_X1 port map( A1 => w(0), A2 => n5, B1 => x(0), B2 => n6, ZN => 
                           n70);
   U98 : NOR2_X1 port map( A1 => n84, A2 => sel(1), ZN => n6);
   U99 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n5);
   U100 : AOI22_X1 port map( A1 => y(0), A2 => n77, B1 => z(0), B2 => n74, ZN 
                           => n69);
   U101 : NOR2_X1 port map( A1 => n85, A2 => n84, ZN => n8);
   U102 : NOR2_X1 port map( A1 => n85, A2 => sel(0), ZN => n7);
   U103 : CLKBUF_X1 port map( A => n8, Z => n74);
   U110 : CLKBUF_X1 port map( A => n5, Z => n83);
   U111 : CLKBUF_X1 port map( A => n7, Z => n77);
   U112 : CLKBUF_X1 port map( A => n6, Z => n80);
   U113 : INV_X1 port map( A => sel(1), ZN => n85);
   U114 : INV_X1 port map( A => sel(0), ZN => n84);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity sign_ext_alt_N_IN016_N_IN18_N_OUT32 is

   port( ctrl_in, zero_padding : in std_logic;  data_in : in std_logic_vector 
         (15 downto 0);  data_ext : out std_logic_vector (31 downto 0));

end sign_ext_alt_N_IN016_N_IN18_N_OUT32;

architecture SYN_dflow of sign_ext_alt_N_IN016_N_IN18_N_OUT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal data_ext_30_port, data_ext_15_port, data_ext_14_port, 
      data_ext_13_port, data_ext_12_port, data_ext_11_port, data_ext_10_port, 
      data_ext_9_port, data_ext_8_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, data_ext_31_port, n15, n16 : std_logic;

begin
   data_ext <= ( data_ext_31_port, data_ext_30_port, data_ext_31_port, 
      data_ext_30_port, data_ext_31_port, data_ext_30_port, data_ext_31_port, 
      data_ext_30_port, data_ext_31_port, data_ext_30_port, data_ext_31_port, 
      data_ext_30_port, data_ext_31_port, data_ext_30_port, data_ext_31_port, 
      data_ext_31_port, data_ext_15_port, data_ext_14_port, data_ext_13_port, 
      data_ext_12_port, data_ext_11_port, data_ext_10_port, data_ext_9_port, 
      data_ext_8_port, data_in(7), data_in(6), data_in(5), data_in(4), 
      data_in(3), data_in(2), data_in(1), data_in(0) );
   
   U4 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => data_ext_9_port);
   U5 : NAND2_X1 port map( A1 => data_in(9), A2 => ctrl_in, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n5, ZN => data_ext_8_port);
   U7 : NAND2_X1 port map( A1 => data_in(8), A2 => ctrl_in, ZN => n5);
   U8 : OAI21_X1 port map( B1 => n16, B2 => n6, A => n3, ZN => data_ext_30_port
                           );
   U9 : OR2_X1 port map( A1 => n15, A2 => zero_padding, ZN => n6);
   U10 : OAI21_X1 port map( B1 => n15, B2 => n16, A => n3, ZN => 
                           data_ext_15_port);
   U11 : NAND2_X1 port map( A1 => n3, A2 => n7, ZN => data_ext_14_port);
   U12 : NAND2_X1 port map( A1 => data_in(14), A2 => ctrl_in, ZN => n7);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n8, ZN => data_ext_13_port);
   U14 : NAND2_X1 port map( A1 => data_in(13), A2 => ctrl_in, ZN => n8);
   U15 : NAND2_X1 port map( A1 => n3, A2 => n9, ZN => data_ext_12_port);
   U16 : NAND2_X1 port map( A1 => data_in(12), A2 => ctrl_in, ZN => n9);
   U17 : NAND2_X1 port map( A1 => n3, A2 => n10, ZN => data_ext_11_port);
   U18 : NAND2_X1 port map( A1 => data_in(11), A2 => ctrl_in, ZN => n10);
   U19 : NAND2_X1 port map( A1 => n3, A2 => n11, ZN => data_ext_10_port);
   U20 : NAND2_X1 port map( A1 => data_in(10), A2 => ctrl_in, ZN => n11);
   U21 : NAND2_X1 port map( A1 => n12, A2 => data_in(7), ZN => n3);
   U22 : NOR2_X1 port map( A1 => zero_padding, A2 => ctrl_in, ZN => n12);
   U3 : CLKBUF_X1 port map( A => data_ext_30_port, Z => data_ext_31_port);
   U23 : INV_X1 port map( A => ctrl_in, ZN => n15);
   U24 : INV_X1 port map( A => data_in(15), ZN => n16);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_3 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_3;

architecture SYN_behav of gen_reg_N32_3 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n107, n116, n117, n118, n119, n120, n121, n122, n123,
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n171, B2 => n107, A => n147, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n107, A2 => data_in(23), ZN => n147);
   U4 : OAI21_X1 port map( B1 => n172, B2 => n97, A => n146, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n107, ZN => n146);
   U6 : OAI21_X1 port map( B1 => n173, B2 => ld, A => n145, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => n97, ZN => n145);
   U8 : OAI21_X1 port map( B1 => n174, B2 => n98, A => n144, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => n97, ZN => n144);
   U10 : OAI21_X1 port map( B1 => n175, B2 => ld, A => n143, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => n107, ZN => n143);
   U12 : OAI21_X1 port map( B1 => n176, B2 => n107, A => n142, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => n107, ZN => n142);
   U14 : OAI21_X1 port map( B1 => n148, B2 => n97, A => n141, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => n107, ZN => n141);
   U16 : OAI21_X1 port map( B1 => n149, B2 => ld, A => n140, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n107, ZN => n140);
   U18 : OAI21_X1 port map( B1 => n150, B2 => n97, A => n139, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n107, ZN => n139);
   U20 : OAI21_X1 port map( B1 => n177, B2 => n97, A => n138, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n107, ZN => n138);
   U22 : OAI21_X1 port map( B1 => n151, B2 => n98, A => n137, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n107, ZN => n137);
   U24 : OAI21_X1 port map( B1 => n152, B2 => n107, A => n136, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n107, ZN => n136);
   U26 : OAI21_X1 port map( B1 => n153, B2 => n107, A => n135, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n107, ZN => n135);
   U28 : OAI21_X1 port map( B1 => n154, B2 => n98, A => n134, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n107, ZN => n134);
   U30 : OAI21_X1 port map( B1 => n155, B2 => n97, A => n133, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n107, ZN => n133);
   U32 : OAI21_X1 port map( B1 => n156, B2 => n98, A => n132, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n107, ZN => n132);
   U34 : OAI21_X1 port map( B1 => n157, B2 => n107, A => n131, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n107, ZN => n131);
   U36 : OAI21_X1 port map( B1 => n158, B2 => n97, A => n130, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n98, ZN => n130);
   U38 : OAI21_X1 port map( B1 => n159, B2 => n98, A => n129, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n107, ZN => n129);
   U40 : OAI21_X1 port map( B1 => n160, B2 => n98, A => n128, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n97, ZN => n128);
   U42 : OAI21_X1 port map( B1 => n178, B2 => n98, A => n127, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => n98, ZN => n127);
   U44 : OAI21_X1 port map( B1 => n161, B2 => n97, A => n126, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n97, ZN => n126);
   U46 : OAI21_X1 port map( B1 => n162, B2 => n107, A => n125, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => n98, ZN => n125);
   U48 : OAI21_X1 port map( B1 => n163, B2 => n98, A => n124, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n97, ZN => n124);
   U50 : OAI21_X1 port map( B1 => n164, B2 => ld, A => n123, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n98, ZN => n123);
   U52 : OAI21_X1 port map( B1 => n165, B2 => n98, A => n122, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n97, ZN => n122);
   U54 : OAI21_X1 port map( B1 => n166, B2 => n97, A => n121, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n98, ZN => n121);
   U56 : OAI21_X1 port map( B1 => n167, B2 => n98, A => n120, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n97, ZN => n120);
   U58 : OAI21_X1 port map( B1 => n168, B2 => n97, A => n119, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n119);
   U60 : OAI21_X1 port map( B1 => n169, B2 => n97, A => n118, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n97, ZN => n118);
   U62 : OAI21_X1 port map( B1 => n170, B2 => n107, A => n117, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n117);
   U64 : OAI21_X1 port map( B1 => n179, B2 => n98, A => n116, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n107, ZN => n116);
   U70 : CLKBUF_X1 port map( A => n107, Z => n97);
   U71 : CLKBUF_X1 port map( A => n107, Z => n98);
   U79 : CLKBUF_X1 port map( A => ld, Z => n107);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n179);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n178);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n177);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n176);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n175);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n174);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n173);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n172);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n171);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n170);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n169);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n168);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n167);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n166);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n165);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n164);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n163);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n162);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n161);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n160);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n159);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n158);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n157);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n156);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n155);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n154);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n153);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n152);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n151);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n150);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n149);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n148);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_mux21_N32_1 is

   port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m : 
         out std_logic_vector (31 downto 0));

end gen_mux21_N32_1;

architecture SYN_dflow of gen_mux21_N32_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n68, n70 : std_logic;

begin
   
   U34 : AOI22_X1 port map( A1 => x(9), A2 => n33, B1 => y(9), B2 => n68, ZN =>
                           n34);
   U35 : AOI22_X1 port map( A1 => x(8), A2 => n33, B1 => y(8), B2 => sel, ZN =>
                           n35);
   U36 : AOI22_X1 port map( A1 => x(7), A2 => n70, B1 => y(7), B2 => n68, ZN =>
                           n36);
   U37 : AOI22_X1 port map( A1 => x(6), A2 => n33, B1 => y(6), B2 => n68, ZN =>
                           n37);
   U38 : AOI22_X1 port map( A1 => x(5), A2 => n33, B1 => y(5), B2 => sel, ZN =>
                           n38);
   U39 : AOI22_X1 port map( A1 => x(4), A2 => n33, B1 => y(4), B2 => n68, ZN =>
                           n39);
   U40 : AOI22_X1 port map( A1 => x(3), A2 => n70, B1 => y(3), B2 => n68, ZN =>
                           n40);
   U41 : AOI22_X1 port map( A1 => x(31), A2 => n33, B1 => y(31), B2 => sel, ZN 
                           => n41);
   U42 : AOI22_X1 port map( A1 => x(30), A2 => n70, B1 => y(30), B2 => n68, ZN 
                           => n42);
   U43 : AOI22_X1 port map( A1 => x(2), A2 => n33, B1 => y(2), B2 => sel, ZN =>
                           n43);
   U44 : AOI22_X1 port map( A1 => x(29), A2 => n70, B1 => y(29), B2 => n68, ZN 
                           => n44);
   U45 : AOI22_X1 port map( A1 => x(28), A2 => n33, B1 => y(28), B2 => sel, ZN 
                           => n45);
   U46 : AOI22_X1 port map( A1 => x(27), A2 => n70, B1 => y(27), B2 => sel, ZN 
                           => n46);
   U47 : AOI22_X1 port map( A1 => x(26), A2 => n70, B1 => y(26), B2 => n68, ZN 
                           => n47);
   U48 : AOI22_X1 port map( A1 => x(25), A2 => n70, B1 => y(25), B2 => sel, ZN 
                           => n48);
   U49 : AOI22_X1 port map( A1 => x(24), A2 => n70, B1 => y(24), B2 => n68, ZN 
                           => n49);
   U50 : AOI22_X1 port map( A1 => x(23), A2 => n70, B1 => y(23), B2 => n68, ZN 
                           => n50);
   U51 : AOI22_X1 port map( A1 => x(22), A2 => n70, B1 => y(22), B2 => n68, ZN 
                           => n51);
   U52 : AOI22_X1 port map( A1 => x(21), A2 => n70, B1 => y(21), B2 => n68, ZN 
                           => n52);
   U53 : AOI22_X1 port map( A1 => x(20), A2 => n70, B1 => y(20), B2 => n68, ZN 
                           => n53);
   U54 : AOI22_X1 port map( A1 => x(1), A2 => n70, B1 => y(1), B2 => n68, ZN =>
                           n54);
   U55 : AOI22_X1 port map( A1 => x(19), A2 => n70, B1 => y(19), B2 => n68, ZN 
                           => n55);
   U56 : AOI22_X1 port map( A1 => x(18), A2 => n70, B1 => y(18), B2 => n68, ZN 
                           => n56);
   U57 : AOI22_X1 port map( A1 => x(17), A2 => n70, B1 => y(17), B2 => n68, ZN 
                           => n57);
   U58 : AOI22_X1 port map( A1 => x(16), A2 => n70, B1 => y(16), B2 => n68, ZN 
                           => n58);
   U59 : AOI22_X1 port map( A1 => x(15), A2 => n70, B1 => y(15), B2 => n68, ZN 
                           => n59);
   U60 : AOI22_X1 port map( A1 => x(14), A2 => n70, B1 => y(14), B2 => n68, ZN 
                           => n60);
   U61 : AOI22_X1 port map( A1 => x(13), A2 => n70, B1 => y(13), B2 => sel, ZN 
                           => n61);
   U62 : AOI22_X1 port map( A1 => x(12), A2 => n70, B1 => y(12), B2 => n68, ZN 
                           => n62);
   U63 : AOI22_X1 port map( A1 => x(11), A2 => n70, B1 => y(11), B2 => sel, ZN 
                           => n63);
   U64 : AOI22_X1 port map( A1 => x(10), A2 => n70, B1 => y(10), B2 => sel, ZN 
                           => n64);
   U65 : AOI22_X1 port map( A1 => x(0), A2 => n70, B1 => y(0), B2 => sel, ZN =>
                           n65);
   U2 : CLKBUF_X1 port map( A => n70, Z => n33);
   U3 : INV_X1 port map( A => sel, ZN => n70);
   U9 : INV_X1 port map( A => n65, ZN => m(0));
   U10 : INV_X1 port map( A => n54, ZN => m(1));
   U11 : INV_X1 port map( A => n43, ZN => m(2));
   U12 : INV_X1 port map( A => n64, ZN => m(10));
   U13 : INV_X1 port map( A => n63, ZN => m(11));
   U14 : INV_X1 port map( A => n62, ZN => m(12));
   U15 : INV_X1 port map( A => n61, ZN => m(13));
   U16 : INV_X1 port map( A => n60, ZN => m(14));
   U17 : INV_X1 port map( A => n59, ZN => m(15));
   U18 : INV_X1 port map( A => n58, ZN => m(16));
   U19 : INV_X1 port map( A => n57, ZN => m(17));
   U20 : INV_X1 port map( A => n56, ZN => m(18));
   U21 : INV_X1 port map( A => n55, ZN => m(19));
   U22 : INV_X1 port map( A => n53, ZN => m(20));
   U23 : INV_X1 port map( A => n52, ZN => m(21));
   U24 : INV_X1 port map( A => n51, ZN => m(22));
   U25 : INV_X1 port map( A => n50, ZN => m(23));
   U26 : INV_X1 port map( A => n49, ZN => m(24));
   U27 : INV_X1 port map( A => n48, ZN => m(25));
   U28 : INV_X1 port map( A => n47, ZN => m(26));
   U29 : INV_X1 port map( A => n46, ZN => m(27));
   U30 : INV_X1 port map( A => n45, ZN => m(28));
   U31 : INV_X1 port map( A => n44, ZN => m(29));
   U32 : INV_X1 port map( A => n42, ZN => m(30));
   U33 : INV_X1 port map( A => n40, ZN => m(3));
   U66 : INV_X1 port map( A => n39, ZN => m(4));
   U67 : INV_X1 port map( A => n38, ZN => m(5));
   U68 : INV_X1 port map( A => n37, ZN => m(6));
   U69 : INV_X1 port map( A => n36, ZN => m(7));
   U70 : INV_X1 port map( A => n35, ZN => m(8));
   U71 : INV_X1 port map( A => n34, ZN => m(9));
   U72 : INV_X1 port map( A => n41, ZN => m(31));
   U74 : CLKBUF_X1 port map( A => sel, Z => n68);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_mux21_N32_2 is

   port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m : 
         out std_logic_vector (31 downto 0));

end gen_mux21_N32_2;

architecture SYN_dflow of gen_mux21_N32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n67, n70 : std_logic;

begin
   
   U34 : AOI22_X1 port map( A1 => x(9), A2 => n70, B1 => y(9), B2 => n67, ZN =>
                           n34);
   U35 : AOI22_X1 port map( A1 => x(8), A2 => n33, B1 => y(8), B2 => n67, ZN =>
                           n35);
   U36 : AOI22_X1 port map( A1 => x(7), A2 => n33, B1 => y(7), B2 => n67, ZN =>
                           n36);
   U37 : AOI22_X1 port map( A1 => x(6), A2 => n33, B1 => y(6), B2 => n67, ZN =>
                           n37);
   U38 : AOI22_X1 port map( A1 => x(5), A2 => n70, B1 => y(5), B2 => n67, ZN =>
                           n38);
   U39 : AOI22_X1 port map( A1 => x(4), A2 => n33, B1 => y(4), B2 => n67, ZN =>
                           n39);
   U40 : AOI22_X1 port map( A1 => x(3), A2 => n70, B1 => y(3), B2 => n67, ZN =>
                           n40);
   U41 : AOI22_X1 port map( A1 => x(31), A2 => n33, B1 => y(31), B2 => sel, ZN 
                           => n41);
   U42 : AOI22_X1 port map( A1 => x(30), A2 => n33, B1 => y(30), B2 => n67, ZN 
                           => n42);
   U43 : AOI22_X1 port map( A1 => x(2), A2 => n33, B1 => y(2), B2 => n67, ZN =>
                           n43);
   U44 : AOI22_X1 port map( A1 => x(29), A2 => n70, B1 => y(29), B2 => n67, ZN 
                           => n44);
   U45 : AOI22_X1 port map( A1 => x(28), A2 => n33, B1 => y(28), B2 => n67, ZN 
                           => n45);
   U46 : AOI22_X1 port map( A1 => x(27), A2 => n70, B1 => y(27), B2 => n67, ZN 
                           => n46);
   U47 : AOI22_X1 port map( A1 => x(26), A2 => n70, B1 => y(26), B2 => n67, ZN 
                           => n47);
   U48 : AOI22_X1 port map( A1 => x(25), A2 => n70, B1 => y(25), B2 => n67, ZN 
                           => n48);
   U49 : AOI22_X1 port map( A1 => x(24), A2 => n70, B1 => y(24), B2 => sel, ZN 
                           => n49);
   U50 : AOI22_X1 port map( A1 => x(23), A2 => n70, B1 => y(23), B2 => n67, ZN 
                           => n50);
   U51 : AOI22_X1 port map( A1 => x(22), A2 => n70, B1 => y(22), B2 => sel, ZN 
                           => n51);
   U52 : AOI22_X1 port map( A1 => x(21), A2 => n70, B1 => y(21), B2 => n67, ZN 
                           => n52);
   U53 : AOI22_X1 port map( A1 => x(20), A2 => n70, B1 => y(20), B2 => n67, ZN 
                           => n53);
   U54 : AOI22_X1 port map( A1 => x(1), A2 => n70, B1 => y(1), B2 => n67, ZN =>
                           n54);
   U55 : AOI22_X1 port map( A1 => x(19), A2 => n70, B1 => y(19), B2 => n67, ZN 
                           => n55);
   U56 : AOI22_X1 port map( A1 => x(18), A2 => n70, B1 => y(18), B2 => n67, ZN 
                           => n56);
   U57 : AOI22_X1 port map( A1 => x(17), A2 => n70, B1 => y(17), B2 => n67, ZN 
                           => n57);
   U58 : AOI22_X1 port map( A1 => x(16), A2 => n70, B1 => y(16), B2 => n67, ZN 
                           => n58);
   U59 : AOI22_X1 port map( A1 => x(15), A2 => n70, B1 => y(15), B2 => sel, ZN 
                           => n59);
   U60 : AOI22_X1 port map( A1 => x(14), A2 => n70, B1 => y(14), B2 => n67, ZN 
                           => n60);
   U61 : AOI22_X1 port map( A1 => x(13), A2 => n70, B1 => y(13), B2 => sel, ZN 
                           => n61);
   U62 : AOI22_X1 port map( A1 => x(12), A2 => n70, B1 => y(12), B2 => sel, ZN 
                           => n62);
   U63 : AOI22_X1 port map( A1 => x(11), A2 => n70, B1 => y(11), B2 => n67, ZN 
                           => n63);
   U64 : AOI22_X1 port map( A1 => x(10), A2 => n70, B1 => y(10), B2 => n67, ZN 
                           => n64);
   U65 : AOI22_X1 port map( A1 => x(0), A2 => n70, B1 => y(0), B2 => n67, ZN =>
                           n65);
   U2 : CLKBUF_X1 port map( A => n70, Z => n33);
   U3 : INV_X1 port map( A => sel, ZN => n70);
   U9 : INV_X1 port map( A => n40, ZN => m(3));
   U10 : INV_X1 port map( A => n39, ZN => m(4));
   U11 : INV_X1 port map( A => n37, ZN => m(6));
   U12 : INV_X1 port map( A => n36, ZN => m(7));
   U13 : INV_X1 port map( A => n54, ZN => m(1));
   U14 : INV_X1 port map( A => n43, ZN => m(2));
   U15 : INV_X1 port map( A => n38, ZN => m(5));
   U16 : INV_X1 port map( A => n35, ZN => m(8));
   U17 : INV_X1 port map( A => n34, ZN => m(9));
   U18 : INV_X1 port map( A => n57, ZN => m(17));
   U19 : INV_X1 port map( A => n56, ZN => m(18));
   U20 : INV_X1 port map( A => n55, ZN => m(19));
   U21 : INV_X1 port map( A => n53, ZN => m(20));
   U22 : INV_X1 port map( A => n52, ZN => m(21));
   U23 : INV_X1 port map( A => n48, ZN => m(25));
   U24 : INV_X1 port map( A => n47, ZN => m(26));
   U25 : INV_X1 port map( A => n46, ZN => m(27));
   U26 : INV_X1 port map( A => n45, ZN => m(28));
   U27 : INV_X1 port map( A => n44, ZN => m(29));
   U28 : INV_X1 port map( A => n42, ZN => m(30));
   U29 : INV_X1 port map( A => n51, ZN => m(22));
   U30 : INV_X1 port map( A => n50, ZN => m(23));
   U31 : INV_X1 port map( A => n49, ZN => m(24));
   U32 : INV_X1 port map( A => n41, ZN => m(31));
   U33 : CLKBUF_X1 port map( A => sel, Z => n67);
   U66 : INV_X1 port map( A => n65, ZN => m(0));
   U67 : INV_X1 port map( A => n64, ZN => m(10));
   U68 : INV_X1 port map( A => n63, ZN => m(11));
   U69 : INV_X1 port map( A => n62, ZN => m(12));
   U70 : INV_X1 port map( A => n61, ZN => m(13));
   U71 : INV_X1 port map( A => n60, ZN => m(14));
   U72 : INV_X1 port map( A => n59, ZN => m(15));
   U73 : INV_X1 port map( A => n58, ZN => m(16));

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity cpsr is

   port( clk, rst, ld, FL3, FL2, FL1, FL0 : in std_logic;  N, Z, C, V : out 
         std_logic);

end cpsr;

architecture SYN_status of cpsr is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal Z_port, n9, n10, n1, n2, n4, n5, net83865, n6, n7, n11, n12, n14, n15
      , n_1064 : std_logic;

begin
   Z <= Z_port;
   
   U2 : OAI21_X1 port map( B1 => n4, B2 => ld, A => n5, ZN => n9);
   U3 : NAND2_X1 port map( A1 => ld, A2 => FL1, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n7, A2 => net83865, ZN => n6);
   U7 : NAND2_X1 port map( A1 => FL0, A2 => ld, ZN => n7);
   U9 : NAND2_X1 port map( A1 => n12, A2 => n14, ZN => n11);
   U10 : NAND2_X1 port map( A1 => FL3, A2 => ld, ZN => n12);
   U12 : OR2_X1 port map( A1 => n2, A2 => ld, ZN => n14);
   U13 : OR2_X1 port map( A1 => n1, A2 => ld, ZN => net83865);
   Z_reg : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => Z_port, QN =>
                           n_1064);
   C_reg : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => C, QN => n4);
   V_reg : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => V, QN => n1);
   N_reg : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => N, QN => n2);
   U4 : INV_X1 port map( A => ld, ZN => n15);
   U5 : MUX2_X1 port map( A => FL2, B => Z_port, S => n15, Z => n10);

end SYN_status;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_5 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_5;

architecture SYN_behav of gen_reg_N32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n34, net75165, net75159, net76910, net76909, net76918, net76917
      , net82841, n97, n98, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n156, B2 => net75165, A => n132, ZN => n9);
   U3 : NAND2_X1 port map( A1 => net76918, A2 => data_in(23), ZN => n132);
   U4 : OAI21_X1 port map( B1 => n157, B2 => net75165, A => n131, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => net76917, ZN => n131);
   U6 : OAI21_X1 port map( B1 => n158, B2 => net76910, A => n130, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => net76917, ZN => n130);
   U8 : OAI21_X1 port map( B1 => n159, B2 => net76909, A => n129, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => net76918, ZN => n129);
   U10 : OAI21_X1 port map( B1 => n160, B2 => net76910, A => n128, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => net76917, ZN => n128);
   U12 : OAI21_X1 port map( B1 => n161, B2 => net75165, A => n127, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => net76917, ZN => n127);
   U14 : OAI21_X1 port map( B1 => n133, B2 => net76910, A => n126, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => net76918, ZN => n126);
   U16 : OAI21_X1 port map( B1 => n134, B2 => net75165, A => n125, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => net76918, ZN => n125);
   U18 : OAI21_X1 port map( B1 => n135, B2 => net75159, A => n124, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => net76918, ZN => n124);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n98, ZN => n123);
   U22 : OAI21_X1 port map( B1 => n136, B2 => net76917, A => n122, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => net76918, ZN => n122);
   U24 : OAI21_X1 port map( B1 => n137, B2 => net76918, A => n121, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n98, ZN => n121);
   U26 : OAI21_X1 port map( B1 => n138, B2 => net75159, A => n120, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => net76918, ZN => n120);
   U28 : OAI21_X1 port map( B1 => n139, B2 => net76918, A => n119, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n98, ZN => n119);
   U30 : OAI21_X1 port map( B1 => n140, B2 => net76917, A => n118, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => net76918, ZN => n118);
   U32 : OAI21_X1 port map( B1 => n141, B2 => net75159, A => n117, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n98, ZN => n117);
   U34 : OAI21_X1 port map( B1 => n142, B2 => n98, A => n116, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => net76918, ZN => n116);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ld, A => n115, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n98, ZN => n115);
   U38 : OAI21_X1 port map( B1 => n144, B2 => ld, A => n114, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => net76918, ZN => n114);
   U40 : OAI21_X1 port map( B1 => n145, B2 => net76918, A => n113, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n98, ZN => n113);
   U44 : OAI21_X1 port map( B1 => n146, B2 => net76909, A => n112, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n98, ZN => n112);
   U46 : OAI21_X1 port map( B1 => n147, B2 => net75165, A => n111, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => net76918, ZN => n111);
   U48 : OAI21_X1 port map( B1 => n148, B2 => net76909, A => n110, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n98, ZN => n110);
   U50 : OAI21_X1 port map( B1 => n149, B2 => net76909, A => n109, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => net75165, ZN => n109);
   U52 : OAI21_X1 port map( B1 => n150, B2 => net76910, A => n108, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n98, ZN => n108);
   U54 : OAI21_X1 port map( B1 => n151, B2 => net76910, A => n107, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n98, ZN => n107);
   U56 : OAI21_X1 port map( B1 => n152, B2 => net76910, A => n106, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n98, ZN => n106);
   U58 : OAI21_X1 port map( B1 => n153, B2 => net76909, A => n105, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n105);
   U60 : OAI21_X1 port map( B1 => n154, B2 => net76909, A => n104, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n98, ZN => n104);
   U62 : OAI21_X1 port map( B1 => n155, B2 => net76909, A => n103, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => net75165, ZN => n103);
   U64 : OAI21_X1 port map( B1 => n163, B2 => net76910, A => n102, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n98, ZN => n102);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => net76917, ZN => n97);
   U66 : NAND2_X1 port map( A1 => n97, A2 => net82841, ZN => n2);
   U67 : OR2_X1 port map( A1 => n34, A2 => n98, ZN => net82841);
   U72 : CLKBUF_X1 port map( A => ld, Z => n98);
   U76 : CLKBUF_X1 port map( A => net75159, Z => net76917);
   U77 : CLKBUF_X1 port map( A => ld, Z => net76918);
   U78 : CLKBUF_X1 port map( A => net75165, Z => net76909);
   U79 : CLKBUF_X1 port map( A => net75165, Z => net76910);
   U83 : CLKBUF_X1 port map( A => ld, Z => net75159);
   U85 : CLKBUF_X1 port map( A => ld, Z => net75165);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n34);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n162);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n161);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n160);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n159);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n158);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n157);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n156);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n155);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n154);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n153);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n152);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n151);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n150);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n149);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n148);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n147);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n146);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n145);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n144);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n143);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n142);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n141);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n140);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n139);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n138);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n137);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n136);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n135);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n134);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n133);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n163);
   U20 : OR2_X1 port map( A1 => n162, A2 => net75165, ZN => n164);
   U42 : NAND2_X1 port map( A1 => n123, A2 => n164, ZN => n3);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_N32 is

   port( ALU_OPCODE : in std_logic_vector (0 to 6);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  NEG, ZERO, CARRY, OVF : out std_logic
         ;  OUTALU : out std_logic_vector (31 downto 0));

end ALU_N32;

architecture SYN_ARITH of ALU_N32 is

   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_N32_DW01_addsub_3
      port( A, B : in std_logic_vector (32 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (32 downto 0);  CO : out 
            std_logic);
   end component;
   
   component ALU_N32_DW02_mult_0
      port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_N32_DW01_cmp6_1
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component ALU_N32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N1568, N1572, N1573, N1576, N1577, N1610, N1611, N1612, N1613, N1614,
      N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624, 
      N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, 
      N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1979, N1980, N1981, 
      N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991, 
      N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, 
      N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, 
      U2_U1_Z_0, n1, n2, n3, n4, n259, n260, n261, n262, n263, n264, n265, n266
      , n267, n268, n269, n271, n272, n273, n274, n275, n278, n279, n280, n281,
      n282, n283, n284, n285, n286, n287, n288, n289, n291, n292, n294, n295, 
      n301, n302, n305, n306, n308, n309, n310, n311, n312, n313, n314, n315, 
      n320, n321, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n502, n503, n504, n506, 
      n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n522, 
      n524, n526, n527, n528, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n562, 
      n563, n564, n565, n566, n567, n568, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n623, n624, n625, 
      n626, n627, n628, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n665, n666, n667, n668, n669, n670, n671, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n762, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
      n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, 
      n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, 
      n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, 
      n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, 
      n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
      n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, 
      n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, 
      n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, 
      n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, 
      n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
      n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, 
      n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, 
      n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, 
      n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
      n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
      n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
      n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, 
      n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, 
      n1166, n1167, n1168, n1169, n1170, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1195, n1199, n1200, n1201, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
      n1234, n1235, n1236, n1239, n1240, n1241, n1242, n1243, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1339, net74224, net74225, net74226, net74227, net74229, net74231,
      net74234, net74235, net74236, net74238, net74243, net74247, net74248, 
      net74250, net74252, net74253, net74264, net74284, net74293, net74295, 
      net74362, net74365, net74367, net74386, net74400, net74426, net74436, 
      net74444, net74450, net74455, net74463, net74464, net76217, net76297, 
      net76311, net76329, net76327, net76325, net76555, net76617, net76624, 
      net76732, net77046, net77050, net77055, net82287, net82473, net82699, 
      net82733, net82773, net82835, net82867, net82891, net82890, net82949, 
      net83048, net83091, net83203, net83207, net83238, net83237, net74233, 
      n509, net83853, net83851, net83893, net83926, net83941, net83955, n307, 
      n304, net86262, net83085, n251, n250, net87741, net87738, net87788, 
      net88905, net88934, net88949, net82508, net77056, net77027, n254, n252, 
      n249, n297, net92254, net92255, net92271, net92300, net83880, net82650, 
      n318, n317, net92259, net83925, n303, n300, n299, n298, n296, n362, n630,
      n629, n622, n270, n508, n1238, n1237, net82307, net83927, net82381, 
      net74249, net74228, n505, n1244, net82880, net76321, net86253, net82819, 
      net82639, net74246, net74222, n363, n1338, n1171, n1194, n1196, n1198, 
      n1340, n1341, n1343, n1344, n1345, n1346, n1348, n1349, n1350, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1359, n1361, n1363, n1364, n1365, 
      n1367, n1369, n1370, n1371, n1373, n1376, n1377, n1378, n1381, n1383, 
      n1384, n1385, n1386, n1387, n1391, n1392, n1393, n1394, n1397, n1399, 
      n1401, n1403, n1404, n1405, n1407, n1409, n1414, n1415, n1416, n1418, 
      n1420, n1421, n1422, n1424, n1425, n1426, n1427, n1429, n1430, n1432, 
      n1436, n1437, n1438, n1440, n1447, n1448, n1450, n1452, n1453, n1456, 
      n1457, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1470, n1471, n1472, n1474, n1475, n1481, n1532, n1535, n1538, 
      n1540, n1545, n1549, n1551, n1555, n1561, n1568_port, n1573_port, 
      n1577_port, n1582, n1585, n1588, n1589, n1595, n1597, n1598, n1599, n1600
      , n1601, n1604, n1605, n1606, n1607, n1608, n1609, n1610_port, n1611_port
      , n1612_port, n1613_port, n1614_port, n1615_port, n1616_port, n1617_port,
      n1618_port, n1619_port, n1620_port, n1621_port, n1622_port, n1624_port, 
      n1625_port, n1626_port, n1627_port, n1628_port, n1629_port, n1630_port, 
      n1631_port, n1632_port, n1633_port, n1634_port, n1635_port, n1636_port, 
      n1637_port, n1638_port, n1639_port, n1640_port, n1641_port, n1642, n1643,
      n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, 
      n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, 
      n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, 
      n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
      n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
      n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, 
      n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, 
      n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
      n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, 
      n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
      n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1797, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   n3 <= '1';
   n4 <= '0';
   U259 : NOR4_X1 port map( A1 => net74450, A2 => n261, A3 => n262, A4 => n263,
                           ZN => n260);
   U260 : NOR4_X1 port map( A1 => n265, A2 => n266, A3 => n267, A4 => n268, ZN 
                           => n259);
   U265 : NOR4_X1 port map( A1 => n1609, A2 => n1608, A3 => n279, A4 => n280, 
                           ZN => n278);
   U270 : NOR4_X1 port map( A1 => n1598, A2 => n1597, A3 => n291, A4 => 
                           net74444, ZN => n286);
   U282 : NOR2_X1 port map( A1 => n311, A2 => net74238, ZN => n309);
   U283 : OAI21_X1 port map( B1 => n312, B2 => net83091, A => n313, ZN => n305)
                           ;
   U284 : AOI22_X1 port map( A1 => net92254, A2 => net74226, B1 => n314, B2 => 
                           net74238, ZN => n312);
   U285 : NAND2_X1 port map( A1 => n315, A2 => net83085, ZN => n295);
   U293 : OAI21_X1 port map( B1 => n324, B2 => net76321, A => n325, ZN => 
                           OUTALU(9));
   U294 : NAND2_X1 port map( A1 => n291, A2 => net74246, ZN => n325);
   U295 : OAI21_X1 port map( B1 => n281, B2 => net76321, A => n326, ZN => 
                           OUTALU(8));
   U296 : NAND2_X1 port map( A1 => n1609, A2 => net74246, ZN => n326);
   U297 : NOR4_X1 port map( A1 => n327, A2 => n328, A3 => n329, A4 => n330, ZN 
                           => n324);
   U298 : AOI21_X1 port map( B1 => n331, B2 => n1653, A => n1618_port, ZN => 
                           n330);
   U299 : OAI21_X1 port map( B1 => n1713, B2 => n333, A => n334, ZN => n332);
   U300 : AOI22_X1 port map( A1 => n1655, A2 => n335, B1 => n1656, B2 => n336, 
                           ZN => n334);
   U301 : AOI21_X1 port map( B1 => n337, B2 => n1657, A => n338, ZN => n331);
   U302 : OAI21_X1 port map( B1 => n1658, B2 => n339, A => n1660, ZN => n338);
   U303 : AOI21_X1 port map( B1 => n340, B2 => n1386, A => n1650, ZN => n329);
   U304 : AOI22_X1 port map( A1 => DATA1(9), A2 => net76217, B1 => n1385, B2 =>
                           n1758, ZN => n340);
   U305 : OAI21_X1 port map( B1 => n1726, B2 => n1668, A => n342, ZN => n328);
   U306 : AOI21_X1 port map( B1 => DATA1(9), B2 => n343, A => n344, ZN => n342)
                           ;
   U307 : OAI21_X1 port map( B1 => n1416, B2 => n345, A => net76311, ZN => n343
                           );
   U308 : NAND2_X1 port map( A1 => n347, A2 => n348, ZN => n327);
   U309 : AOI22_X1 port map( A1 => n349, A2 => n350, B1 => n351, B2 => net82287
                           , ZN => n348);
   U310 : OR2_X1 port map( A1 => n353, A2 => n354, ZN => n349);
   U311 : OAI21_X1 port map( B1 => n1713, B2 => n1675, A => n355, ZN => n354);
   U312 : AOI22_X1 port map( A1 => n1549, A2 => n335, B1 => n357, B2 => n336, 
                           ZN => n355);
   U313 : OAI21_X1 port map( B1 => n1715, B2 => n1664, A => n358, ZN => n353);
   U314 : AOI22_X1 port map( A1 => n359, A2 => n360, B1 => n361, B2 => n337, ZN
                           => n358);
   U315 : AOI22_X1 port map( A1 => N1619, A2 => net76325, B1 => N1988, B2 => 
                           n362, ZN => n347);
   U316 : OAI21_X1 port map( B1 => net76617, B2 => n281, A => n364, ZN => 
                           OUTALU(7));
   U317 : NAND2_X1 port map( A1 => net76617, A2 => n279, ZN => n364);
   U318 : NOR4_X1 port map( A1 => n365, A2 => n366, A3 => n367, A4 => n368, ZN 
                           => n281);
   U319 : NAND2_X1 port map( A1 => n369, A2 => n370, ZN => n368);
   U320 : AOI22_X1 port map( A1 => N1618, A2 => net76325, B1 => N1987, B2 => 
                           n362, ZN => n369);
   U321 : OAI21_X1 port map( B1 => net74362, B2 => n371, A => n372, ZN => n367)
                           ;
   U322 : AOI22_X1 port map( A1 => n373, A2 => n374, B1 => n375, B2 => n376, ZN
                           => n372);
   U323 : OAI21_X1 port map( B1 => n1707, B2 => n377, A => n378, ZN => n366);
   U324 : AOI22_X1 port map( A1 => n1460, A2 => n379, B1 => n380, B2 => n381, 
                           ZN => n378);
   U325 : NAND2_X1 port map( A1 => n382, A2 => net76311, ZN => n379);
   U326 : AOI22_X1 port map( A1 => DATA1(8), A2 => n341, B1 => net76297, B2 => 
                           n1759, ZN => n382);
   U327 : OAI21_X1 port map( B1 => n383, B2 => n1665, A => n384, ZN => n365);
   U328 : AOI21_X1 port map( B1 => DATA1(8), B2 => n385, A => n386, ZN => n384)
                           ;
   U329 : NOR3_X1 port map( A1 => n1658, A2 => n387, A3 => n1618_port, ZN => 
                           n386);
   U330 : OAI21_X1 port map( B1 => n1460, B2 => n345, A => n1386, ZN => n385);
   U331 : OAI21_X1 port map( B1 => n1607, B2 => net76321, A => n389, ZN => 
                           OUTALU(6));
   U332 : NAND2_X1 port map( A1 => n279, A2 => net74246, ZN => n389);
   U334 : OAI21_X1 port map( B1 => n394, B2 => n1716, A => n395, ZN => n393);
   U335 : AOI21_X1 port map( B1 => n396, B2 => DATA1(7), A => n344, ZN => n395)
                           ;
   U336 : OAI21_X1 port map( B1 => n345, B2 => n1457, A => net76311, ZN => n396
                           );
   U337 : AOI22_X1 port map( A1 => n397, A2 => n398, B1 => n399, B2 => n350, ZN
                           => n392);
   U338 : NAND2_X1 port map( A1 => n400, A2 => n401, ZN => n399);
   U339 : AOI21_X1 port map( B1 => n361, B2 => n402, A => n403, ZN => n401);
   U340 : OAI21_X1 port map( B1 => n1687, B2 => net74367, A => n404, ZN => n403
                           );
   U341 : NAND2_X1 port map( A1 => n405, A2 => n406, ZN => n404);
   U342 : AOI22_X1 port map( A1 => n356, A2 => n408, B1 => n357, B2 => n409, ZN
                           => n400);
   U343 : AOI22_X1 port map( A1 => n1457, A2 => n410, B1 => n411, B2 => n412, 
                           ZN => n391);
   U344 : OR2_X1 port map( A1 => n413, A2 => n414, ZN => n412);
   U345 : OAI21_X1 port map( B1 => n1719, B2 => n415, A => n416, ZN => n414);
   U346 : AOI22_X1 port map( A1 => n1657, A2 => n402, B1 => n1655, B2 => n408, 
                           ZN => n416);
   U347 : OAI21_X1 port map( B1 => n1678, B2 => n1658, A => n417, ZN => n413);
   U348 : AOI21_X1 port map( B1 => n1652, B2 => n406, A => n418, ZN => n417);
   U349 : NAND2_X1 port map( A1 => n420, A2 => net76311, ZN => n410);
   U350 : AOI22_X1 port map( A1 => DATA1(7), A2 => n341, B1 => net76297, B2 => 
                           n1760, ZN => n420);
   U351 : AOI22_X1 port map( A1 => N1617, A2 => net76325, B1 => N1986, B2 => 
                           n362, ZN => n390);
   U352 : OAI21_X1 port map( B1 => n285, B2 => net76321, A => n421, ZN => 
                           OUTALU(5));
   U353 : NAND2_X1 port map( A1 => n280, A2 => net74246, ZN => n421);
   U355 : OAI21_X1 port map( B1 => n394, B2 => n1731, A => n426, ZN => n425);
   U356 : AOI21_X1 port map( B1 => n427, B2 => DATA1(6), A => n344, ZN => n426)
                           ;
   U358 : AOI22_X1 port map( A1 => n397, A2 => n428, B1 => n429, B2 => n350, ZN
                           => n424);
   U359 : NAND2_X1 port map( A1 => n430, A2 => n431, ZN => n429);
   U360 : AOI21_X1 port map( B1 => n361, B2 => n432, A => n433, ZN => n431);
   U361 : OAI21_X1 port map( B1 => n1686, B2 => net74367, A => n434, ZN => n433
                           );
   U362 : NAND2_X1 port map( A1 => n405, A2 => n435, ZN => n434);
   U363 : AOI22_X1 port map( A1 => n356, A2 => n437, B1 => n1545, B2 => n438, 
                           ZN => n430);
   U364 : AOI22_X1 port map( A1 => net82473, A2 => n439, B1 => n411, B2 => n440
                           , ZN => n423);
   U365 : OR2_X1 port map( A1 => n441, A2 => n442, ZN => n440);
   U366 : OAI21_X1 port map( B1 => n1723, B2 => n415, A => n443, ZN => n442);
   U367 : AOI22_X1 port map( A1 => n1657, A2 => n432, B1 => n1655, B2 => n437, 
                           ZN => n443);
   U368 : OAI21_X1 port map( B1 => n1729, B2 => n333, A => n444, ZN => n441);
   U369 : AOI21_X1 port map( B1 => n445, B2 => n446, A => n418, ZN => n444);
   U370 : NAND2_X1 port map( A1 => n447, A2 => net76311, ZN => n439);
   U371 : AOI22_X1 port map( A1 => DATA1(6), A2 => n341, B1 => net76297, B2 => 
                           n1761, ZN => n447);
   U372 : AOI22_X1 port map( A1 => N1616, A2 => net76325, B1 => N1985, B2 => 
                           n362, ZN => n422);
   U373 : OAI21_X1 port map( B1 => net76617, B2 => n285, A => n448, ZN => 
                           OUTALU(4));
   U374 : NAND2_X1 port map( A1 => net76617, A2 => n282, ZN => n448);
   U375 : NOR3_X1 port map( A1 => n449, A2 => n450, A3 => n451, ZN => n285);
   U376 : OAI21_X1 port map( B1 => n1727, B2 => n1668, A => n452, ZN => n451);
   U377 : OAI21_X1 port map( B1 => n453, B2 => n454, A => n350, ZN => n452);
   U378 : OAI21_X1 port map( B1 => n1713, B2 => n1672, A => n455, ZN => n454);
   U379 : AOI22_X1 port map( A1 => n357, A2 => n335, B1 => n456, B2 => n336, ZN
                           => n455);
   U380 : NAND2_X1 port map( A1 => n457, A2 => n458, ZN => n453);
   U381 : AOI22_X1 port map( A1 => n459, A2 => net76732, B1 => n359, B2 => n460
                           , ZN => n458);
   U382 : NOR2_X1 port map( A1 => n1714, A2 => n1688, ZN => n459);
   U383 : AOI22_X1 port map( A1 => n1549, A2 => n337, B1 => n405, B2 => n461, 
                           ZN => n457);
   U384 : OAI21_X1 port map( B1 => n462, B2 => n394, A => n463, ZN => n450);
   U385 : AOI21_X1 port map( B1 => DATA1(5), B2 => n464, A => n344, ZN => n463)
                           ;
   U386 : OAI21_X1 port map( B1 => n1456, B2 => n345, A => net76311, ZN => n464
                           );
   U387 : NAND2_X1 port map( A1 => n1532, A2 => net82287, ZN => n394);
   U388 : NAND2_X1 port map( A1 => n466, A2 => n467, ZN => n449);
   U389 : AOI22_X1 port map( A1 => n1456, A2 => n468, B1 => n411, B2 => n469, 
                           ZN => n467);
   U390 : NAND2_X1 port map( A1 => n470, A2 => n471, ZN => n469);
   U391 : AOI21_X1 port map( B1 => n461, B2 => n1652, A => n1654, ZN => n471);
   U392 : AOI22_X1 port map( A1 => n1655, A2 => n337, B1 => n1656, B2 => n335, 
                           ZN => n472);
   U393 : AOI21_X1 port map( B1 => n473, B2 => n1657, A => n474, ZN => n470);
   U394 : OAI21_X1 port map( B1 => n1658, B2 => n475, A => n1660, ZN => n474);
   U395 : NAND2_X1 port map( A1 => n476, A2 => n1386, ZN => n468);
   U396 : AOI22_X1 port map( A1 => DATA1(5), A2 => n341, B1 => n1385, B2 => 
                           n1762, ZN => n476);
   U397 : AOI22_X1 port map( A1 => N1615, A2 => net76325, B1 => N1984, B2 => 
                           n362, ZN => n466);
   U398 : OAI21_X1 port map( B1 => n1605, B2 => net76321, A => n477, ZN => 
                           OUTALU(3));
   U399 : NAND2_X1 port map( A1 => n282, A2 => net74246, ZN => n477);
   U401 : NOR3_X1 port map( A1 => n482, A2 => n483, A3 => n484, ZN => n481);
   U402 : OAI33_X1 port map( A1 => n485, A2 => n1403, A3 => net74362, B1 => 
                           n1658, B2 => n486, B3 => n1618_port, ZN => n484);
   U403 : NOR2_X1 port map( A1 => n487, A2 => n1763, ZN => n483);
   U404 : AOI21_X1 port map( B1 => n1385, B2 => net74367, A => net76555, ZN => 
                           n487);
   U405 : OAI21_X1 port map( B1 => n1708, B2 => n377, A => n489, ZN => n482);
   U406 : AOI22_X1 port map( A1 => net76732, A2 => n490, B1 => n380, B2 => n491
                           , ZN => n489);
   U407 : OAI21_X1 port map( B1 => n1618_port, B2 => n492, A => n493, ZN => 
                           n380);
   U408 : NAND2_X1 port map( A1 => n356, A2 => n350, ZN => n493);
   U409 : NAND2_X1 port map( A1 => n494, A2 => n495, ZN => n490);
   U410 : AOI22_X1 port map( A1 => n1685, A2 => n350, B1 => DATA1(4), B2 => 
                           net76217, ZN => n495);
   U411 : AOI21_X1 port map( B1 => n1385, B2 => n1763, A => net76555, ZN => 
                           n494);
   U412 : AOI21_X1 port map( B1 => n411, B2 => n1657, A => n497, ZN => n377);
   U413 : NOR2_X1 port map( A1 => n1672, A2 => net74247, ZN => n497);
   U414 : AOI21_X1 port map( B1 => N1983, B2 => n362, A => n1614_port, ZN => 
                           n480);
   U415 : AOI21_X1 port map( B1 => n418, B2 => n411, A => n344, ZN => n370);
   U416 : NAND2_X1 port map( A1 => N1614, A2 => net76327, ZN => n479);
   U417 : AOI22_X1 port map( A1 => n373, A2 => n381, B1 => n375, B2 => n498, ZN
                           => n478);
   U418 : OAI21_X1 port map( B1 => n333, B2 => n1618_port, A => n1674, ZN => 
                           n375);
   U419 : OAI21_X1 port map( B1 => n1618_port, B2 => n415, A => n499, ZN => 
                           n373);
   U420 : NAND2_X1 port map( A1 => n1545, A2 => n350, ZN => n499);
   U421 : OAI21_X1 port map( B1 => net77055, B2 => net76321, A => n1775, ZN => 
                           OUTALU(31));
   U428 : OAI21_X1 port map( B1 => n510, B2 => n1646, A => n511, ZN => n504);
   U429 : AOI22_X1 port map( A1 => n1555, A2 => n513, B1 => n514, B2 => n515, 
                           ZN => n511);
   U430 : NAND2_X1 port map( A1 => n516, A2 => n517, ZN => n515);
   U431 : AOI21_X1 port map( B1 => DATA1(30), B2 => n518, A => n519, ZN => n517
                           );
   U432 : AOI22_X1 port map( A1 => n1573_port, A2 => DATA1(28), B1 => 
                           n1568_port, B2 => DATA1(29), ZN => n516);
   U436 : OAI21_X1 port map( B1 => n302, B2 => n528, A => net92271, ZN => n527)
                           ;
   U437 : NAND2_X1 port map( A1 => n531, A2 => n532, ZN => n502);
   U438 : AOI22_X1 port map( A1 => DATA1(31), A2 => n533, B1 => n534, B2 => 
                           n1735, ZN => n532);
   U439 : OAI21_X1 port map( B1 => DATA2(31), B2 => n345, A => net76311, ZN => 
                           n533);
   U440 : AOI22_X1 port map( A1 => n1666, A2 => n535, B1 => DATA2(31), B2 => 
                           n536, ZN => n531);
   U441 : NAND2_X1 port map( A1 => n537, A2 => net76311, ZN => n536);
   U442 : AOI22_X1 port map( A1 => DATA1(31), A2 => n341, B1 => n1385, B2 => 
                           net74284, ZN => n537);
   U443 : OAI21_X1 port map( B1 => n1601, B2 => net76321, A => n538, ZN => 
                           OUTALU(2));
   U444 : NAND2_X1 port map( A1 => n283, A2 => net74246, ZN => n538);
   U446 : NOR3_X1 port map( A1 => n543, A2 => n544, A3 => n545, ZN => n542);
   U447 : NOR3_X1 port map( A1 => n546, A2 => n547, A3 => net74367, ZN => n545)
                           ;
   U448 : NOR2_X1 port map( A1 => n548, A2 => n1764, ZN => n543);
   U449 : AOI21_X1 port map( B1 => n1385, B2 => n1692, A => net76555, ZN => 
                           n548);
   U450 : AOI21_X1 port map( B1 => n388, B2 => n1683, A => n549, ZN => n541);
   U451 : AOI21_X1 port map( B1 => n550, B2 => n551, A => n552, ZN => n549);
   U452 : AOI21_X1 port map( B1 => n1532, B2 => n406, A => n553, ZN => n551);
   U453 : NOR2_X1 port map( A1 => n554, A2 => n1693, ZN => n553);
   U454 : NOR4_X1 port map( A1 => n555, A2 => n556, A3 => n557, A4 => n558, ZN 
                           => n554);
   U455 : NOR2_X1 port map( A1 => n1577_port, A2 => n1762, ZN => n558);
   U456 : NAND2_X1 port map( A1 => n559, A2 => n560, ZN => n406);
   U457 : AOI22_X1 port map( A1 => DATA1(7), A2 => n1582, B1 => DATA1(6), B2 =>
                           n1475, ZN => n560);
   U458 : AOI22_X1 port map( A1 => DATA1(9), A2 => n1573_port, B1 => DATA1(8), 
                           B2 => n1481, ZN => n559);
   U459 : AOI22_X1 port map( A1 => n1540, A2 => n402, B1 => n1538, B2 => n408, 
                           ZN => n550);
   U460 : AOI22_X1 port map( A1 => n1403, A2 => n565, B1 => n1551, B2 => n566, 
                           ZN => n540);
   U461 : NAND2_X1 port map( A1 => n567, A2 => net76311, ZN => n565);
   U462 : AOI22_X1 port map( A1 => n1404, A2 => n341, B1 => n1385, B2 => n1764,
                           ZN => n567);
   U463 : AOI22_X1 port map( A1 => N1613, A2 => net76327, B1 => N1982, B2 => 
                           n362, ZN => n539);
   U464 : OAI21_X1 port map( B1 => n1604, B2 => net76321, A => n568, ZN => 
                           OUTALU(29));
   U465 : NAND2_X1 port map( A1 => n284, A2 => net74246, ZN => n568);
   U467 : AOI21_X1 port map( B1 => DATA1(30), B2 => n573, A => n574, ZN => n572
                           );
   U468 : OAI21_X1 port map( B1 => n1621_port, B2 => n575, A => n1610_port, ZN 
                           => n574);
   U469 : NAND2_X1 port map( A1 => n1535, A2 => n577, ZN => n575);
   U470 : OAI21_X1 port map( B1 => DATA2(30), B2 => n345, A => net76311, ZN => 
                           n573);
   U471 : AOI22_X1 port map( A1 => n534, A2 => n578, B1 => DATA2(30), B2 => 
                           n579, ZN => n571);
   U472 : NAND2_X1 port map( A1 => n580, A2 => net76311, ZN => n579);
   U473 : AOI22_X1 port map( A1 => DATA1(30), A2 => net76217, B1 => n1385, B2 
                           => n1740, ZN => n580);
   U474 : AOI22_X1 port map( A1 => n581, A2 => n582, B1 => n1438, B2 => n1768, 
                           ZN => n570);
   U475 : NAND2_X1 port map( A1 => n583, A2 => n584, ZN => n581);
   U476 : NOR3_X1 port map( A1 => n585, A2 => n586, A3 => n587, ZN => n584);
   U478 : AOI21_X1 port map( B1 => n589, B2 => n590, A => n1675, ZN => n586);
   U479 : AOI21_X1 port map( B1 => DATA1(29), B2 => n1582, A => n591, ZN => 
                           n590);
   U480 : AOI22_X1 port map( A1 => DATA1(27), A2 => n520, B1 => n1481, B2 => 
                           DATA1(28), ZN => n589);
   U482 : AOI22_X1 port map( A1 => n357, A2 => n593, B1 => net76732, B2 => n594
                           , ZN => n583);
   U484 : OAI21_X1 port map( B1 => net74436, B2 => net76321, A => n595, ZN => 
                           OUTALU(28));
   U485 : NAND2_X1 port map( A1 => n1429, A2 => net74246, ZN => n595);
   U487 : AOI21_X1 port map( B1 => n600, B2 => n360, A => n601, ZN => n599);
   U488 : OAI21_X1 port map( B1 => n1693, B2 => n1621_port, A => n1674, ZN => 
                           n600);
   U489 : NOR2_X1 port map( A1 => n1675, A2 => net74247, ZN => n534);
   U490 : AOI22_X1 port map( A1 => DATA1(29), A2 => n602, B1 => DATA2(29), B2 
                           => n603, ZN => n598);
   U491 : NAND2_X1 port map( A1 => n604, A2 => net76311, ZN => n603);
   U492 : AOI22_X1 port map( A1 => DATA1(29), A2 => net76217, B1 => n1385, B2 
                           => n1741, ZN => n604);
   U493 : OAI21_X1 port map( B1 => DATA2(29), B2 => n345, A => net76311, ZN => 
                           n602);
   U494 : AOI22_X1 port map( A1 => n605, A2 => n582, B1 => n1448, B2 => n1768, 
                           ZN => n597);
   U495 : OR2_X1 port map( A1 => n606, A2 => n607, ZN => n605);
   U496 : OAI21_X1 port map( B1 => n1725, B2 => n1664, A => n608, ZN => n607);
   U497 : AOI22_X1 port map( A1 => n356, A2 => n609, B1 => n357, B2 => n610, ZN
                           => n608);
   U498 : NAND2_X1 port map( A1 => n612, A2 => n613, ZN => n606);
   U499 : AOI21_X1 port map( B1 => net76732, B2 => n614, A => n615, ZN => n613)
                           ;
   U500 : AOI21_X1 port map( B1 => n616, B2 => n617, A => n1675, ZN => n615);
   U501 : AOI22_X1 port map( A1 => DATA1(28), A2 => n518, B1 => n1561, B2 => 
                           DATA1(29), ZN => n617);
   U502 : AOI22_X1 port map( A1 => DATA1(26), A2 => n520, B1 => DATA1(27), B2 
                           => n1568_port, ZN => n616);
   U503 : AOI22_X1 port map( A1 => n359, A2 => n346, B1 => n361, B2 => n618, ZN
                           => n612);
   U505 : AOI22_X1 port map( A1 => n272, A2 => net74246, B1 => n273, B2 => 
                           net76617, ZN => n619);
   U507 : AOI21_X1 port map( B1 => DATA1(28), B2 => n624, A => n625, ZN => n623
                           );
   U508 : OAI21_X1 port map( B1 => n1693, B2 => n626, A => n1610_port, ZN => 
                           n625);
   U509 : NOR2_X1 port map( A1 => net74426, A2 => net74248, ZN => n601);
   U510 : OR2_X1 port map( A1 => n1704, A2 => n627, ZN => n626);
   U511 : OAI21_X1 port map( B1 => DATA2(28), B2 => n345, A => net76311, ZN => 
                           n624);
   U515 : AOI22_X1 port map( A1 => n631, A2 => n582, B1 => net83048, B2 => 
                           n1768, ZN => n621);
   U516 : OR2_X1 port map( A1 => n632, A2 => n633, ZN => n631);
   U517 : OAI21_X1 port map( B1 => n1712, B2 => n1672, A => n634, ZN => n633);
   U518 : AOI22_X1 port map( A1 => n1545, A2 => n635, B1 => n456, B2 => n636, 
                           ZN => n634);
   U519 : NAND2_X1 port map( A1 => n637, A2 => n638, ZN => n632);
   U520 : AOI21_X1 port map( B1 => n359, B2 => n639, A => n640, ZN => n638);
   U521 : NOR3_X1 port map( A1 => n485, A2 => n1692, A3 => net74367, ZN => n640
                           );
   U522 : AOI22_X1 port map( A1 => n405, A2 => n641, B1 => n1549, B2 => n642, 
                           ZN => n637);
   U523 : AOI22_X1 port map( A1 => N1638, A2 => net76327, B1 => N2007, B2 => 
                           n362, ZN => n620);
   U524 : AOI22_X1 port map( A1 => n273, A2 => net74246, B1 => net76617, B2 => 
                           n274, ZN => n643);
   U526 : NOR4_X1 port map( A1 => n648, A2 => n649, A3 => n650, A4 => n651, ZN 
                           => n647);
   U527 : NOR3_X1 port map( A1 => n1667, A2 => n1718, A3 => n1693, ZN => n651);
   U528 : OAI21_X1 port map( B1 => n652, B2 => net74365, A => n653, ZN => n649)
                           ;
   U529 : OAI21_X1 port map( B1 => n654, B2 => net76555, A => DATA1(27), ZN => 
                           n653);
   U530 : NOR2_X1 port map( A1 => DATA2(27), A2 => n345, ZN => n654);
   U531 : NAND2_X1 port map( A1 => n655, A2 => n656, ZN => n648);
   U532 : AOI22_X1 port map( A1 => n1666, A2 => n657, B1 => n658, B2 => n659, 
                           ZN => n656);
   U533 : AOI22_X1 port map( A1 => DATA2(27), A2 => n660, B1 => n661, B2 => 
                           n662, ZN => n655);
   U534 : NAND2_X1 port map( A1 => n663, A2 => n1386, ZN => n660);
   U535 : AOI22_X1 port map( A1 => DATA1(27), A2 => n341, B1 => n1385, B2 => 
                           n1742, ZN => n663);
   U538 : NAND2_X1 port map( A1 => N1637, A2 => net76327, ZN => n665);
   U539 : AOI22_X1 port map( A1 => n1671, A2 => n666, B1 => n1670, B2 => n524, 
                           ZN => n645);
   U540 : AOI22_X1 port map( A1 => n1555, A2 => n530, B1 => n514, B2 => n513, 
                           ZN => n644);
   U541 : NAND2_X1 port map( A1 => n667, A2 => n668, ZN => n513);
   U542 : AOI22_X1 port map( A1 => DATA1(26), A2 => n1582, B1 => DATA1(27), B2 
                           => n1561, ZN => n668);
   U543 : AOI22_X1 port map( A1 => DATA1(24), A2 => n1573_port, B1 => DATA1(25)
                           , B2 => n1481, ZN => n667);
   U544 : OAI21_X1 port map( B1 => n1355, B2 => net76321, A => n669, ZN => 
                           OUTALU(25));
   U545 : NAND2_X1 port map( A1 => n274, A2 => net74246, ZN => n669);
   U547 : NOR4_X1 port map( A1 => n674, A2 => n675, A3 => n650, A4 => n676, ZN 
                           => n673);
   U548 : NOR3_X1 port map( A1 => n1667, A2 => n1722, A3 => n1693, ZN => n676);
   U549 : OAI21_X1 port map( B1 => n1732, B2 => net74365, A => n677, ZN => n675
                           );
   U550 : OAI21_X1 port map( B1 => n678, B2 => net76555, A => DATA1(26), ZN => 
                           n677);
   U551 : NOR2_X1 port map( A1 => DATA2(26), A2 => n345, ZN => n678);
   U552 : NOR2_X1 port map( A1 => n1667, A2 => n1696, ZN => n628);
   U553 : NAND2_X1 port map( A1 => n679, A2 => n680, ZN => n674);
   U554 : AOI22_X1 port map( A1 => n1666, A2 => n681, B1 => n658, B2 => n682, 
                           ZN => n680);
   U555 : AOI22_X1 port map( A1 => DATA2(26), A2 => n683, B1 => n661, B2 => 
                           n1689, ZN => n679);
   U556 : NAND2_X1 port map( A1 => n685, A2 => net76311, ZN => n683);
   U557 : AOI22_X1 port map( A1 => DATA1(26), A2 => n341, B1 => n1385, B2 => 
                           n1743, ZN => n685);
   U560 : NAND2_X1 port map( A1 => N1636, A2 => net76327, ZN => n687);
   U561 : AOI22_X1 port map( A1 => n1671, A2 => n688, B1 => n1670, B2 => n593, 
                           ZN => n671);
   U562 : AOI22_X1 port map( A1 => n1555, A2 => n592, B1 => n1551, B2 => n588, 
                           ZN => n670);
   U563 : NAND2_X1 port map( A1 => n689, A2 => n690, ZN => n588);
   U564 : AOI21_X1 port map( B1 => DATA1(25), B2 => n1582, A => n691, ZN => 
                           n690);
   U565 : AOI22_X1 port map( A1 => DATA1(26), A2 => n1561, B1 => DATA1(24), B2 
                           => n1568_port, ZN => n689);
   U566 : OAI21_X1 port map( B1 => net76617, B2 => n1355, A => n692, ZN => 
                           OUTALU(24));
   U567 : NAND2_X1 port map( A1 => net76617, A2 => n1381, ZN => n692);
   U570 : AOI22_X1 port map( A1 => n1416, A2 => n1768, B1 => N1635, B2 => 
                           net76327, ZN => n697);
   U571 : NAND2_X1 port map( A1 => n698, A2 => n699, ZN => n695);
   U572 : AOI22_X1 port map( A1 => n1671, A2 => n611, B1 => n1670, B2 => n610, 
                           ZN => n699);
   U573 : AOI22_X1 port map( A1 => n1555, A2 => n609, B1 => n514, B2 => n618, 
                           ZN => n698);
   U574 : NAND2_X1 port map( A1 => n700, A2 => n701, ZN => n618);
   U575 : AOI22_X1 port map( A1 => DATA1(24), A2 => n1582, B1 => DATA1(25), B2 
                           => n1561, ZN => n701);
   U576 : AOI22_X1 port map( A1 => DATA1(22), A2 => n1573_port, B1 => DATA1(23)
                           , B2 => n1481, ZN => n700);
   U577 : OAI21_X1 port map( B1 => n339, B2 => n1621_port, A => n702, ZN => 
                           n694);
   U578 : AOI22_X1 port map( A1 => n703, A2 => n704, B1 => DATA2(25), B2 => 
                           n705, ZN => n702);
   U579 : NAND2_X1 port map( A1 => n706, A2 => n1386, ZN => n705);
   U580 : AOI22_X1 port map( A1 => DATA1(25), A2 => net76217, B1 => n1385, B2 
                           => n1744, ZN => n706);
   U581 : NOR2_X1 port map( A1 => n704, A2 => n707, ZN => n339);
   U582 : OAI21_X1 port map( B1 => n1714, B2 => n1696, A => n708, ZN => n704);
   U583 : NAND2_X1 port map( A1 => n576, A2 => n460, ZN => n708);
   U584 : NAND2_X1 port map( A1 => n709, A2 => n710, ZN => n693);
   U585 : AOI21_X1 port map( B1 => DATA1(25), B2 => n711, A => n650, ZN => n710
                           );
   U586 : OAI21_X1 port map( B1 => DATA2(25), B2 => n345, A => net76311, ZN => 
                           n711);
   U587 : AOI22_X1 port map( A1 => n1666, A2 => n351, B1 => n658, B2 => n346, 
                           ZN => n709);
   U588 : OAI21_X1 port map( B1 => n1727, B2 => n1696, A => n712, ZN => n351);
   U589 : NAND2_X1 port map( A1 => n1540, A2 => n1736, ZN => n712);
   U590 : OAI21_X1 port map( B1 => n714, B2 => net76321, A => n715, ZN => 
                           OUTALU(23));
   U591 : NAND2_X1 port map( A1 => n1381, A2 => net74246, ZN => n715);
   U592 : NAND2_X1 port map( A1 => n716, A2 => n717, ZN => n275);
   U593 : NOR4_X1 port map( A1 => n718, A2 => n719, A3 => n720, A4 => n721, ZN 
                           => n717);
   U594 : AOI21_X1 port map( B1 => n722, B2 => n1386, A => n1628_port, ZN => 
                           n721);
   U595 : AOI22_X1 port map( A1 => DATA1(24), A2 => net76217, B1 => net76297, 
                           B2 => n1745, ZN => n722);
   U596 : NOR2_X1 port map( A1 => n371, A2 => n713, ZN => n720);
   U597 : AOI21_X1 port map( B1 => n1540, B2 => n723, A => n1695, ZN => n371);
   U598 : AOI22_X1 port map( A1 => n576, A2 => n639, B1 => n1532, B2 => n725, 
                           ZN => n724);
   U599 : OAI21_X1 port map( B1 => n726, B2 => n1745, A => n1611_port, ZN => 
                           n719);
   U600 : AOI21_X1 port map( B1 => n1385, B2 => n1628_port, A => net76555, ZN 
                           => n726);
   U601 : OAI21_X1 port map( B1 => n1699, B2 => n522, A => n727, ZN => n718);
   U602 : AOI22_X1 port map( A1 => n661, A2 => n1691, B1 => n1671, B2 => n636, 
                           ZN => n727);
   U603 : NOR2_X1 port map( A1 => n728, A2 => n707, ZN => n387);
   U606 : AOI22_X1 port map( A1 => n1460, A2 => n1768, B1 => N1634, B2 => 
                           net76329, ZN => n731);
   U607 : OAI21_X1 port map( B1 => n383, B2 => n1667, A => n732, ZN => n729);
   U608 : AOI22_X1 port map( A1 => n1555, A2 => n642, B1 => n1551, B2 => n733, 
                           ZN => n732);
   U609 : AOI21_X1 port map( B1 => n1540, B2 => n519, A => n728, ZN => n383);
   U610 : OAI21_X1 port map( B1 => n1704, B2 => n1696, A => n734, ZN => n728);
   U611 : NAND2_X1 port map( A1 => n1535, A2 => n735, ZN => n734);
   U612 : OAI21_X1 port map( B1 => n736, B2 => net76321, A => n737, ZN => 
                           OUTALU(22));
   U613 : NAND2_X1 port map( A1 => n1595, A2 => net74246, ZN => n737);
   U614 : NOR4_X1 port map( A1 => n738, A2 => n739, A3 => n740, A4 => n741, ZN 
                           => n714);
   U615 : OAI21_X1 port map( B1 => net83207, B2 => n1631_port, A => n742, ZN =>
                           n741);
   U616 : AOI22_X1 port map( A1 => n1457, A2 => n1768, B1 => N1633, B2 => 
                           net76329, ZN => n742);
   U617 : NAND2_X1 port map( A1 => n743, A2 => n744, ZN => n740);
   U618 : AOI22_X1 port map( A1 => n1670, A2 => n666, B1 => n1555, B2 => n524, 
                           ZN => n744);
   U619 : AOI22_X1 port map( A1 => n1551, A2 => n530, B1 => n703, B2 => n407, 
                           ZN => n743);
   U620 : OAI21_X1 port map( B1 => n652, B2 => n1688, A => n1694, ZN => n407);
   U621 : NAND2_X1 port map( A1 => n745, A2 => n746, ZN => n530);
   U622 : AOI22_X1 port map( A1 => DATA1(22), A2 => n518, B1 => DATA1(23), B2 
                           => n1475, ZN => n746);
   U623 : AOI22_X1 port map( A1 => DATA1(20), A2 => n1573_port, B1 => DATA1(21)
                           , B2 => n1568_port, ZN => n745);
   U624 : OAI21_X1 port map( B1 => n1720, B2 => n747, A => n748, ZN => n739);
   U625 : AOI22_X1 port map( A1 => DATA2(23), A2 => n749, B1 => n661, B2 => 
                           n419, ZN => n748);
   U626 : NAND2_X1 port map( A1 => n750, A2 => n1694, ZN => n419);
   U627 : OAI21_X1 port map( B1 => n1718, B2 => n1696, A => n752, ZN => n751);
   U628 : NAND2_X1 port map( A1 => n576, A2 => n753, ZN => n752);
   U629 : AOI21_X1 port map( B1 => n1540, B2 => n1734, A => n754, ZN => n750);
   U630 : NAND2_X1 port map( A1 => n755, A2 => n1386, ZN => n749);
   U631 : AOI22_X1 port map( A1 => DATA1(23), A2 => net76217, B1 => n1385, B2 
                           => n1746, ZN => n755);
   U632 : NAND2_X1 port map( A1 => n756, A2 => n757, ZN => n738);
   U633 : AOI21_X1 port map( B1 => DATA1(23), B2 => n758, A => n650, ZN => n757
                           );
   U634 : OAI21_X1 port map( B1 => DATA2(23), B2 => n345, A => net76311, ZN => 
                           n758);
   U635 : AOI22_X1 port map( A1 => n759, A2 => n566, B1 => n658, B2 => n398, ZN
                           => n756);
   U636 : OAI21_X1 port map( B1 => n264, B2 => net76321, A => n760, ZN => 
                           OUTALU(21));
   U637 : NAND2_X1 port map( A1 => n1359, A2 => net74246, ZN => n760);
   U639 : OAI21_X1 port map( B1 => net83207, B2 => n1632_port, A => n765, ZN =>
                           n764);
   U640 : AOI22_X1 port map( A1 => net82473, A2 => n1768, B1 => N1632, B2 => 
                           net76329, ZN => n765);
   U642 : AOI22_X1 port map( A1 => n1670, A2 => n688, B1 => n1555, B2 => n593, 
                           ZN => n767);
   U643 : AOI22_X1 port map( A1 => n514, A2 => n592, B1 => n703, B2 => n436, ZN
                           => n766);
   U644 : OAI21_X1 port map( B1 => n1732, B2 => n1688, A => n768, ZN => n436);
   U645 : NAND2_X1 port map( A1 => n769, A2 => n770, ZN => n592);
   U646 : AOI22_X1 port map( A1 => DATA1(21), A2 => n1582, B1 => DATA1(22), B2 
                           => n1561, ZN => n770);
   U647 : AOI22_X1 port map( A1 => DATA1(19), A2 => n1573_port, B1 => DATA1(20)
                           , B2 => n1481, ZN => n769);
   U648 : OAI21_X1 port map( B1 => n1724, B2 => n747, A => n771, ZN => n762);
   U649 : AOI22_X1 port map( A1 => DATA2(22), A2 => n772, B1 => n661, B2 => 
                           n446, ZN => n771);
   U650 : NAND2_X1 port map( A1 => n773, A2 => n768, ZN => n446);
   U651 : AOI21_X1 port map( B1 => n774, B2 => n1532, A => n775, ZN => n768);
   U653 : AOI21_X1 port map( B1 => n1540, B2 => n577, A => n754, ZN => n773);
   U654 : NAND2_X1 port map( A1 => n777, A2 => n1386, ZN => n772);
   U655 : AOI22_X1 port map( A1 => DATA1(22), A2 => net76217, B1 => net76297, 
                           B2 => n1747, ZN => n777);
   U657 : AOI21_X1 port map( B1 => DATA1(22), B2 => n780, A => n650, ZN => n779
                           );
   U658 : OAI21_X1 port map( B1 => DATA2(22), B2 => n345, A => net76311, ZN => 
                           n780);
   U659 : AOI22_X1 port map( A1 => n759, A2 => n781, B1 => n658, B2 => n428, ZN
                           => n778);
   U661 : NAND2_X1 port map( A1 => net76617, A2 => n262, ZN => n782);
   U663 : OAI21_X1 port map( B1 => net83207, B2 => n1633_port, A => n787, ZN =>
                           n786);
   U664 : AOI22_X1 port map( A1 => n1456, A2 => n1768, B1 => N1631, B2 => 
                           net76329, ZN => n787);
   U665 : NAND2_X1 port map( A1 => n788, A2 => n789, ZN => n785);
   U666 : AOI22_X1 port map( A1 => n1671, A2 => n346, B1 => n1670, B2 => n611, 
                           ZN => n789);
   U667 : AOI22_X1 port map( A1 => n1555, A2 => n610, B1 => n1551, B2 => n609, 
                           ZN => n788);
   U668 : NAND2_X1 port map( A1 => n790, A2 => n791, ZN => n609);
   U669 : AOI22_X1 port map( A1 => DATA1(20), A2 => n1582, B1 => DATA1(21), B2 
                           => n1475, ZN => n791);
   U670 : AOI22_X1 port map( A1 => DATA1(18), A2 => n1573_port, B1 => DATA1(19)
                           , B2 => n1568_port, ZN => n790);
   U671 : OAI21_X1 port map( B1 => n475, B2 => n1621_port, A => n792, ZN => 
                           n784);
   U672 : AOI22_X1 port map( A1 => n703, A2 => n793, B1 => DATA2(21), B2 => 
                           n794, ZN => n792);
   U673 : NAND2_X1 port map( A1 => n795, A2 => n1386, ZN => n794);
   U674 : AOI22_X1 port map( A1 => DATA1(21), A2 => n341, B1 => n1385, B2 => 
                           n1748, ZN => n795);
   U675 : NOR2_X1 port map( A1 => n793, A2 => n754, ZN => n475);
   U676 : OAI21_X1 port map( B1 => n1700, B2 => n1693, A => n796, ZN => n793);
   U677 : AOI22_X1 port map( A1 => n1540, A2 => n360, B1 => n1532, B2 => n460, 
                           ZN => n796);
   U678 : NAND2_X1 port map( A1 => n797, A2 => n798, ZN => n783);
   U679 : AOI21_X1 port map( B1 => DATA1(21), B2 => n799, A => n650, ZN => n798
                           );
   U680 : OAI21_X1 port map( B1 => DATA2(21), B2 => n345, A => n1386, ZN => 
                           n799);
   U681 : AOI22_X1 port map( A1 => n759, A2 => n1736, B1 => n658, B2 => n800, 
                           ZN => n797);
   U682 : NOR2_X1 port map( A1 => n1662, A2 => net74250, ZN => n759);
   U683 : AOI22_X1 port map( A1 => n261, A2 => net74246, B1 => net76617, B2 => 
                           n268, ZN => n801);
   U685 : NOR3_X1 port map( A1 => n806, A2 => n544, A3 => n807, ZN => n805);
   U686 : NOR3_X1 port map( A1 => n546, A2 => n808, A3 => net74367, ZN => n807)
                           ;
   U687 : NOR2_X1 port map( A1 => n809, A2 => n1765, ZN => n806);
   U688 : AOI21_X1 port map( B1 => n1385, B2 => n1698, A => net76555, ZN => 
                           n809);
   U689 : AOI21_X1 port map( B1 => n388, B2 => n1681, A => n810, ZN => n804);
   U690 : AOI21_X1 port map( B1 => n811, B2 => n812, A => n552, ZN => n810);
   U691 : AOI21_X1 port map( B1 => net74367, B2 => n1622_port, A => n703, ZN =>
                           n552);
   U692 : AOI22_X1 port map( A1 => n1535, A2 => n813, B1 => n1532, B2 => n435, 
                           ZN => n812);
   U693 : NAND2_X1 port map( A1 => n814, A2 => n815, ZN => n435);
   U694 : AOI22_X1 port map( A1 => DATA1(6), A2 => n1582, B1 => DATA1(5), B2 =>
                           n1475, ZN => n815);
   U695 : AOI22_X1 port map( A1 => DATA1(8), A2 => n1573_port, B1 => DATA1(7), 
                           B2 => n1481, ZN => n814);
   U696 : NAND2_X1 port map( A1 => n816, A2 => n817, ZN => n813);
   U697 : AOI21_X1 port map( B1 => n1461, B2 => n1582, A => n818, ZN => n817);
   U698 : AOI22_X1 port map( A1 => DATA1(4), A2 => n1573_port, B1 => n1404, B2 
                           => n1568_port, ZN => n816);
   U699 : AOI22_X1 port map( A1 => n1540, A2 => n432, B1 => n1538, B2 => n437, 
                           ZN => n811);
   U700 : NOR2_X1 port map( A1 => net74367, A2 => net74247, ZN => n388);
   U701 : AOI22_X1 port map( A1 => DATA2(2), A2 => n820, B1 => n1551, B2 => 
                           n781, ZN => n803);
   U702 : NAND2_X1 port map( A1 => n821, A2 => n1386, ZN => n820);
   U703 : AOI22_X1 port map( A1 => n1461, A2 => net76217, B1 => net76297, B2 =>
                           n1765, ZN => n821);
   U704 : AOI22_X1 port map( A1 => N1612, A2 => net76325, B1 => N1981, B2 => 
                           n362, ZN => n802);
   U705 : AOI22_X1 port map( A1 => n262, A2 => net74246, B1 => net76617, B2 => 
                           n263, ZN => n822);
   U706 : NAND2_X1 port map( A1 => n823, A2 => n824, ZN => n262);
   U707 : NOR4_X1 port map( A1 => n825, A2 => n1635_port, A3 => n650, A4 => 
                           n826, ZN => n824);
   U708 : NOR3_X1 port map( A1 => n713, A2 => n1403, A3 => n485, ZN => n826);
   U709 : NAND2_X1 port map( A1 => net76732, A2 => n582, ZN => n713);
   U710 : AOI21_X1 port map( B1 => n828, B2 => DATA1(20), A => net74400, ZN => 
                           n827);
   U712 : OAI21_X1 port map( B1 => DATA1(20), B2 => n345, A => n831, ZN => n830
                           );
   U713 : NAND2_X1 port map( A1 => DATA1(20), A2 => net76217, ZN => n831);
   U715 : OAI21_X1 port map( B1 => n1709, B2 => n522, A => n832, ZN => n825);
   U716 : AOI22_X1 port map( A1 => n661, A2 => n1677, B1 => n1671, B2 => n639, 
                           ZN => n832);
   U717 : NOR2_X1 port map( A1 => n833, A2 => n754, ZN => n486);
   U718 : NOR2_X1 port map( A1 => n1679, A2 => net74284, ZN => n754);
   U719 : NOR2_X1 port map( A1 => n834, A2 => n835, ZN => n823);
   U720 : OAI21_X1 port map( B1 => net83207, B2 => n1634_port, A => n836, ZN =>
                           n835);
   U721 : AOI22_X1 port map( A1 => n1768, A2 => net76732, B1 => N1630, B2 => 
                           net76329, ZN => n836);
   U722 : OAI21_X1 port map( B1 => n496, B2 => n1667, A => n837, ZN => n834);
   U723 : AOI22_X1 port map( A1 => n1555, A2 => n635, B1 => n514, B2 => n642, 
                           ZN => n837);
   U724 : AOI21_X1 port map( B1 => n1538, B2 => n519, A => n833, ZN => n496);
   U725 : OAI21_X1 port map( B1 => n1705, B2 => n1696, A => n838, ZN => n833);
   U726 : AOI22_X1 port map( A1 => n1540, A2 => n839, B1 => n1535, B2 => n374, 
                           ZN => n838);
   U727 : AOI22_X1 port map( A1 => n263, A2 => net74246, B1 => net76617, B2 => 
                           n265, ZN => n840);
   U728 : NAND2_X1 port map( A1 => n841, A2 => n842, ZN => n263);
   U729 : NOR4_X1 port map( A1 => n843, A2 => n844, A3 => n845, A4 => n846, ZN 
                           => n842);
   U730 : AOI21_X1 port map( B1 => n847, B2 => n1386, A => n1638_port, ZN => 
                           n846);
   U731 : AOI22_X1 port map( A1 => DATA1(19), A2 => net76217, B1 => n1385, B2 
                           => n1749, ZN => n847);
   U732 : NOR2_X1 port map( A1 => n1716, A2 => n1663, ZN => n845);
   U733 : OAI21_X1 port map( B1 => n848, B2 => n1749, A => n1611_port, ZN => 
                           n844);
   U734 : AOI21_X1 port map( B1 => n1385, B2 => n1638_port, A => net76555, ZN 
                           => n848);
   U735 : OAI21_X1 port map( B1 => n1720, B2 => n522, A => n849, ZN => n843);
   U736 : AOI22_X1 port map( A1 => n661, A2 => n1684, B1 => n1671, B2 => n398, 
                           ZN => n849);
   U737 : AOI21_X1 port map( B1 => n1734, B2 => n1538, A => n850, ZN => n547);
   U738 : NOR2_X1 port map( A1 => n851, A2 => n852, ZN => n841);
   U739 : OAI21_X1 port map( B1 => net83207, B2 => n1636_port, A => n853, ZN =>
                           n852);
   U740 : AOI22_X1 port map( A1 => n1768, A2 => n1403, B1 => N1629, B2 => 
                           net76329, ZN => n853);
   U741 : OAI21_X1 port map( B1 => n564, B2 => n1667, A => n854, ZN => n851);
   U742 : AOI22_X1 port map( A1 => n1555, A2 => n666, B1 => n1551, B2 => n524, 
                           ZN => n854);
   U743 : NAND2_X1 port map( A1 => n855, A2 => n856, ZN => n524);
   U744 : AOI22_X1 port map( A1 => DATA1(18), A2 => n1582, B1 => DATA1(19), B2 
                           => n1475, ZN => n856);
   U745 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1573_port, B1 => DATA1(17)
                           , B2 => n1481, ZN => n855);
   U746 : AOI21_X1 port map( B1 => n1735, B2 => n1538, A => n850, ZN => n564);
   U747 : OAI21_X1 port map( B1 => n1718, B2 => n1688, A => n857, ZN => n850);
   U748 : AOI22_X1 port map( A1 => n576, A2 => n409, B1 => n1532, B2 => n753, 
                           ZN => n857);
   U749 : AOI22_X1 port map( A1 => n265, A2 => net74246, B1 => net76617, B2 => 
                           n266, ZN => n858);
   U750 : NAND2_X1 port map( A1 => n859, A2 => n860, ZN => n265);
   U751 : NOR4_X1 port map( A1 => n861, A2 => n862, A3 => n863, A4 => n864, ZN 
                           => n860);
   U752 : AOI21_X1 port map( B1 => n865, B2 => n1386, A => n1640_port, ZN => 
                           n864);
   U753 : AOI22_X1 port map( A1 => DATA1(18), A2 => net76217, B1 => net76297, 
                           B2 => n1750, ZN => n865);
   U754 : NOR2_X1 port map( A1 => n1731, A2 => n1663, ZN => n863);
   U755 : OAI21_X1 port map( B1 => n866, B2 => n1750, A => n1611_port, ZN => 
                           n862);
   U756 : AOI21_X1 port map( B1 => n1385, B2 => n1640_port, A => net76555, ZN 
                           => n866);
   U757 : OAI21_X1 port map( B1 => n1724, B2 => n522, A => n867, ZN => n861);
   U758 : AOI22_X1 port map( A1 => n661, A2 => n1682, B1 => n1671, B2 => n428, 
                           ZN => n867);
   U759 : AOI21_X1 port map( B1 => n577, B2 => n1538, A => n868, ZN => n808);
   U760 : NOR2_X1 port map( A1 => n869, A2 => n870, ZN => n859);
   U761 : OAI21_X1 port map( B1 => net83207, B2 => n1639_port, A => n871, ZN =>
                           n870);
   U762 : AOI22_X1 port map( A1 => n1768, A2 => DATA2(2), B1 => N1628, B2 => 
                           net76329, ZN => n871);
   U763 : OAI21_X1 port map( B1 => n819, B2 => n1667, A => n872, ZN => n869);
   U764 : AOI22_X1 port map( A1 => n1555, A2 => n688, B1 => n514, B2 => n593, 
                           ZN => n872);
   U765 : NAND2_X1 port map( A1 => n873, A2 => n874, ZN => n593);
   U766 : AOI22_X1 port map( A1 => DATA1(17), A2 => n1582, B1 => DATA1(18), B2 
                           => n1561, ZN => n874);
   U767 : AOI22_X1 port map( A1 => DATA1(15), A2 => n1573_port, B1 => DATA1(16)
                           , B2 => n1481, ZN => n873);
   U768 : AOI21_X1 port map( B1 => n578, B2 => n1538, A => n868, ZN => n819);
   U769 : OAI21_X1 port map( B1 => n1722, B2 => n1688, A => n875, ZN => n868);
   U770 : AOI22_X1 port map( A1 => n1535, A2 => n438, B1 => n1532, B2 => n776, 
                           ZN => n875);
   U771 : AOI22_X1 port map( A1 => n266, A2 => net74246, B1 => net76617, B2 => 
                           n267, ZN => n876);
   U772 : NAND2_X1 port map( A1 => n877, A2 => n878, ZN => n266);
   U773 : NOR4_X1 port map( A1 => n879, A2 => n880, A3 => n881, A4 => n882, ZN 
                           => n878);
   U774 : AOI21_X1 port map( B1 => n883, B2 => n1386, A => n1643, ZN => n882);
   U775 : AOI22_X1 port map( A1 => DATA1(17), A2 => net76217, B1 => net76297, 
                           B2 => n1751, ZN => n883);
   U776 : AOI21_X1 port map( B1 => n884, B2 => n885, A => n627, ZN => n881);
   U777 : AOI22_X1 port map( A1 => n576, A2 => n335, B1 => n1532, B2 => n336, 
                           ZN => n884);
   U778 : NOR2_X1 port map( A1 => n1727, A2 => n747, ZN => n880);
   U779 : OAI21_X1 port map( B1 => n462, B2 => n1663, A => n886, ZN => n879);
   U780 : AOI21_X1 port map( B1 => DATA1(17), B2 => n887, A => n650, ZN => n886
                           );
   U781 : OAI21_X1 port map( B1 => DATA2(17), B2 => n345, A => n1386, ZN => 
                           n887);
   U782 : NOR2_X1 port map( A1 => n888, A2 => n889, ZN => n877);
   U783 : OAI21_X1 port map( B1 => net83207, B2 => n1642, A => n890, ZN => n889
                           );
   U784 : AOI22_X1 port map( A1 => n1768, A2 => DATA2(1), B1 => N1627, B2 => 
                           net76329, ZN => n890);
   U785 : OAI21_X1 port map( B1 => n1728, B2 => n1673, A => n891, ZN => n888);
   U786 : AOI22_X1 port map( A1 => n1670, A2 => n346, B1 => n1555, B2 => n611, 
                           ZN => n891);
   U787 : NAND2_X1 port map( A1 => n892, A2 => n893, ZN => n610);
   U788 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1582, B1 => DATA1(17), B2 
                           => n1561, ZN => n893);
   U789 : AOI22_X1 port map( A1 => DATA1(14), A2 => n1573_port, B1 => DATA1(15)
                           , B2 => n1481, ZN => n892);
   U790 : OAI21_X1 port map( B1 => n894, B2 => net76321, A => n895, ZN => 
                           OUTALU(15));
   U791 : NAND2_X1 port map( A1 => n267, A2 => net74246, ZN => n895);
   U792 : NAND2_X1 port map( A1 => n896, A2 => n897, ZN => n267);
   U793 : NOR4_X1 port map( A1 => n898, A2 => n899, A3 => n900, A4 => n901, ZN 
                           => n897);
   U794 : AOI21_X1 port map( B1 => n902, B2 => n1386, A => n1645, ZN => n901);
   U795 : AOI22_X1 port map( A1 => DATA1(16), A2 => net76217, B1 => n1385, B2 
                           => n1752, ZN => n902);
   U796 : AOI21_X1 port map( B1 => n903, B2 => n1676, A => n627, ZN => n900);
   U797 : NOR2_X1 port map( A1 => n661, A2 => n703, ZN => n627);
   U798 : NOR2_X1 port map( A1 => net74247, A2 => net76732, ZN => n703);
   U799 : NOR2_X1 port map( A1 => n904, A2 => net74248, ZN => n661);
   U800 : AOI22_X1 port map( A1 => n1535, A2 => n381, B1 => n1532, B2 => n374, 
                           ZN => n903);
   U801 : NOR2_X1 port map( A1 => n1711, A2 => n747, ZN => n899);
   U802 : NAND2_X1 port map( A1 => n1545, A2 => n582, ZN => n747);
   U803 : NAND2_X1 port map( A1 => n906, A2 => n907, ZN => n898);
   U804 : AOI21_X1 port map( B1 => n908, B2 => n519, A => n650, ZN => n907);
   U805 : NOR2_X1 port map( A1 => n909, A2 => net74248, ZN => n650);
   U806 : NOR2_X1 port map( A1 => net74247, A2 => n1664, ZN => n908);
   U807 : AOI22_X1 port map( A1 => DATA1(16), A2 => n910, B1 => n658, B2 => 
                           n723, ZN => n906);
   U808 : NOR2_X1 port map( A1 => n1664, A2 => net74250, ZN => n658);
   U809 : OAI21_X1 port map( B1 => DATA2(16), B2 => n345, A => n1386, ZN => 
                           n910);
   U810 : NOR2_X1 port map( A1 => n911, A2 => n912, ZN => n896);
   U811 : OAI21_X1 port map( B1 => net83207, B2 => n1644, A => n913, ZN => n912
                           );
   U812 : AOI22_X1 port map( A1 => n1768, A2 => DATA2(0), B1 => N1626, B2 => 
                           net76327, ZN => n913);
   U813 : OAI21_X1 port map( B1 => n1699, B2 => n1673, A => n914, ZN => n911);
   U814 : AOI22_X1 port map( A1 => n1670, A2 => n639, B1 => n1555, B2 => n636, 
                           ZN => n914);
   U815 : NOR2_X1 port map( A1 => n1672, A2 => net74250, ZN => n512);
   U816 : NAND2_X1 port map( A1 => n1549, A2 => n582, ZN => n522);
   U817 : OAI21_X1 port map( B1 => n915, B2 => net76321, A => n916, ZN => 
                           OUTALU(14));
   U818 : NAND2_X1 port map( A1 => n1600, A2 => net74246, ZN => n916);
   U819 : NOR4_X1 port map( A1 => n917, A2 => n918, A3 => n919, A4 => n920, ZN 
                           => n894);
   U820 : AOI21_X1 port map( B1 => n921, B2 => n1386, A => n1646, ZN => n920);
   U821 : AOI22_X1 port map( A1 => DATA1(15), A2 => net76217, B1 => net76297, 
                           B2 => n1753, ZN => n921);
   U822 : AOI21_X1 port map( B1 => n922, B2 => n923, A => net74247, ZN => n919)
                           ;
   U823 : AOI21_X1 port map( B1 => n361, B2 => n409, A => n924, ZN => n923);
   U824 : OAI21_X1 port map( B1 => n1717, B2 => n1675, A => n925, ZN => n924);
   U825 : NAND2_X1 port map( A1 => n456, A2 => n1735, ZN => n925);
   U826 : AOI22_X1 port map( A1 => n356, A2 => n753, B1 => n357, B2 => n926, ZN
                           => n922);
   U827 : OAI21_X1 port map( B1 => n927, B2 => n1753, A => n1612_port, ZN => 
                           n918);
   U828 : AOI21_X1 port map( B1 => n1385, B2 => n1646, A => net76555, ZN => 
                           n927);
   U829 : NAND2_X1 port map( A1 => n928, A2 => n929, ZN => n917);
   U830 : AOI22_X1 port map( A1 => n411, A2 => n930, B1 => n535, B2 => net82287
                           , ZN => n929);
   U831 : NAND2_X1 port map( A1 => n931, A2 => n932, ZN => n535);
   U832 : AOI22_X1 port map( A1 => n576, A2 => n666, B1 => n1538, B2 => n566, 
                           ZN => n932);
   U833 : NAND2_X1 port map( A1 => n933, A2 => n934, ZN => n666);
   U834 : AOI22_X1 port map( A1 => DATA1(14), A2 => n1582, B1 => DATA1(15), B2 
                           => n1561, ZN => n934);
   U835 : AOI22_X1 port map( A1 => DATA1(12), A2 => n1573_port, B1 => DATA1(13)
                           , B2 => n1481, ZN => n933);
   U836 : AOI22_X1 port map( A1 => n1540, A2 => n398, B1 => n1532, B2 => n659, 
                           ZN => n931);
   U837 : OR2_X1 port map( A1 => n935, A2 => n936, ZN => n930);
   U838 : NAND2_X1 port map( A1 => n937, A2 => n938, ZN => n936);
   U839 : AOI22_X1 port map( A1 => n1655, A2 => n753, B1 => n1656, B2 => n926, 
                           ZN => n937);
   U840 : OAI21_X1 port map( B1 => n1717, B2 => n333, A => n939, ZN => n935);
   U841 : AOI22_X1 port map( A1 => n940, A2 => n1734, B1 => n1657, B2 => n409, 
                           ZN => n939);
   U842 : AOI22_X1 port map( A1 => N1625, A2 => net76325, B1 => N1994, B2 => 
                           n362, ZN => n928);
   U843 : OAI21_X1 port map( B1 => n941, B2 => net76321, A => n942, ZN => 
                           OUTALU(13));
   U844 : NAND2_X1 port map( A1 => n1599, A2 => net74246, ZN => n942);
   U845 : NOR4_X1 port map( A1 => n943, A2 => n944, A3 => n945, A4 => n946, ZN 
                           => n915);
   U846 : AOI21_X1 port map( B1 => n947, B2 => n1386, A => n1647, ZN => n946);
   U847 : AOI22_X1 port map( A1 => DATA1(14), A2 => net76217, B1 => net76297, 
                           B2 => n1754, ZN => n947);
   U848 : AOI21_X1 port map( B1 => n948, B2 => n949, A => net74247, ZN => n945)
                           ;
   U849 : AOI21_X1 port map( B1 => n361, B2 => n438, A => n950, ZN => n949);
   U850 : OAI21_X1 port map( B1 => n1732, B2 => n1664, A => n951, ZN => n950);
   U851 : NAND2_X1 port map( A1 => n405, A2 => n437, ZN => n951);
   U852 : AOI22_X1 port map( A1 => n1549, A2 => n776, B1 => n1545, B2 => n774, 
                           ZN => n948);
   U853 : OAI21_X1 port map( B1 => n952, B2 => n1754, A => n1612_port, ZN => 
                           n944);
   U854 : AOI21_X1 port map( B1 => n1385, B2 => n1647, A => net76555, ZN => 
                           n952);
   U855 : NAND2_X1 port map( A1 => n953, A2 => n954, ZN => n943);
   U856 : AOI22_X1 port map( A1 => n411, A2 => n955, B1 => n594, B2 => net82287
                           , ZN => n954);
   U857 : NAND2_X1 port map( A1 => n956, A2 => n957, ZN => n594);
   U858 : AOI22_X1 port map( A1 => n1535, A2 => n688, B1 => n1538, B2 => n781, 
                           ZN => n957);
   U859 : NAND2_X1 port map( A1 => n958, A2 => n959, ZN => n688);
   U860 : AOI21_X1 port map( B1 => DATA1(13), B2 => n1582, A => n960, ZN => 
                           n959);
   U861 : AOI22_X1 port map( A1 => DATA1(14), A2 => n1475, B1 => DATA1(11), B2 
                           => n1573_port, ZN => n958);
   U862 : AOI22_X1 port map( A1 => n1540, A2 => n428, B1 => n1532, B2 => n682, 
                           ZN => n956);
   U863 : OR2_X1 port map( A1 => n961, A2 => n962, ZN => n955);
   U864 : NAND2_X1 port map( A1 => n963, A2 => n938, ZN => n962);
   U865 : AOI22_X1 port map( A1 => n1655, A2 => n776, B1 => n1656, B2 => n774, 
                           ZN => n963);
   U866 : OAI21_X1 port map( B1 => n1723, B2 => n964, A => n965, ZN => n961);
   U867 : AOI22_X1 port map( A1 => n940, A2 => n577, B1 => n1652, B2 => n437, 
                           ZN => n965);
   U868 : AOI22_X1 port map( A1 => N1624, A2 => net76325, B1 => N1993, B2 => 
                           n362, ZN => n953);
   U869 : OAI21_X1 port map( B1 => n966, B2 => net76321, A => n967, ZN => 
                           OUTALU(12));
   U870 : NAND2_X1 port map( A1 => n1598, A2 => net74246, ZN => n967);
   U871 : NOR4_X1 port map( A1 => n968, A2 => n1613_port, A3 => n969, A4 => 
                           n970, ZN => n941);
   U872 : AOI21_X1 port map( B1 => n971, B2 => n972, A => net74247, ZN => n970)
                           ;
   U873 : AOI21_X1 port map( B1 => n357, B2 => n460, A => n973, ZN => n972);
   U874 : OAI21_X1 port map( B1 => n1714, B2 => n1664, A => n974, ZN => n973);
   U875 : NAND2_X1 port map( A1 => n405, A2 => n337, ZN => n974);
   U876 : AOI22_X1 port map( A1 => n361, A2 => n335, B1 => n356, B2 => n336, ZN
                           => n971);
   U877 : AOI21_X1 port map( B1 => n975, B2 => n1680, A => net74362, ZN => n969
                           );
   U878 : OAI21_X1 port map( B1 => n1727, B2 => n1688, A => n976, ZN => n614);
   U879 : NAND2_X1 port map( A1 => n1538, A2 => n1736, ZN => n976);
   U880 : NAND2_X1 port map( A1 => n977, A2 => n978, ZN => n800);
   U881 : AOI22_X1 port map( A1 => DATA1(4), A2 => n1582, B1 => DATA1(5), B2 =>
                           n1475, ZN => n978);
   U882 : AOI22_X1 port map( A1 => n1461, A2 => n1573_port, B1 => n1404, B2 => 
                           n1481, ZN => n977);
   U883 : AOI22_X1 port map( A1 => n576, A2 => n611, B1 => n1532, B2 => n346, 
                           ZN => n975);
   U884 : NAND2_X1 port map( A1 => n979, A2 => n980, ZN => n346);
   U885 : AOI22_X1 port map( A1 => DATA1(8), A2 => n1582, B1 => DATA1(9), B2 =>
                           n1561, ZN => n980);
   U886 : AOI22_X1 port map( A1 => DATA1(6), A2 => n1573_port, B1 => DATA1(7), 
                           B2 => n1481, ZN => n979);
   U887 : NAND2_X1 port map( A1 => n981, A2 => n982, ZN => n611);
   U888 : AOI22_X1 port map( A1 => DATA1(12), A2 => n1582, B1 => DATA1(13), B2 
                           => n1475, ZN => n982);
   U889 : AOI22_X1 port map( A1 => DATA1(10), A2 => n1573_port, B1 => DATA1(11)
                           , B2 => n1481, ZN => n981);
   U890 : AOI21_X1 port map( B1 => n984, B2 => DATA1(13), A => n344, ZN => n983
                           );
   U891 : OAI21_X1 port map( B1 => n345, B2 => n1448, A => n1386, ZN => n984);
   U892 : NAND2_X1 port map( A1 => n985, A2 => n986, ZN => n968);
   U893 : AOI22_X1 port map( A1 => n1448, A2 => n987, B1 => n411, B2 => n988, 
                           ZN => n986);
   U894 : OR2_X1 port map( A1 => n989, A2 => n990, ZN => n988);
   U895 : NAND2_X1 port map( A1 => n991, A2 => n938, ZN => n990);
   U896 : AOI22_X1 port map( A1 => n1656, A2 => n460, B1 => n1652, B2 => n337, 
                           ZN => n991);
   U897 : OAI21_X1 port map( B1 => n1700, B2 => n492, A => n992, ZN => n989);
   U898 : AOI22_X1 port map( A1 => n940, A2 => n360, B1 => n1657, B2 => n335, 
                           ZN => n992);
   U899 : NAND2_X1 port map( A1 => n993, A2 => net76311, ZN => n987);
   U900 : AOI22_X1 port map( A1 => DATA1(13), A2 => net76217, B1 => net76297, 
                           B2 => n1755, ZN => n993);
   U901 : AOI22_X1 port map( A1 => N1623, A2 => net76325, B1 => N1992, B2 => 
                           n362, ZN => n985);
   U902 : OAI21_X1 port map( B1 => n292, B2 => net76321, A => n994, ZN => 
                           OUTALU(11));
   U903 : NAND2_X1 port map( A1 => n1597, A2 => net74246, ZN => n994);
   U904 : NOR4_X1 port map( A1 => n995, A2 => n996, A3 => n997, A4 => 
                           n1619_port, ZN => n966);
   U905 : OAI21_X1 port map( B1 => n999, B2 => n1000, A => n411, ZN => n998);
   U906 : NAND2_X1 port map( A1 => n1001, A2 => n938, ZN => n1000);
   U907 : AOI21_X1 port map( B1 => n445, B2 => n1002, A => n418, ZN => n938);
   U908 : NOR2_X1 port map( A1 => net74284, A2 => n576, ZN => n1002);
   U909 : AOI22_X1 port map( A1 => n1656, A2 => n735, B1 => n1652, B2 => n491, 
                           ZN => n1001);
   U910 : OAI21_X1 port map( B1 => n1702, B2 => n492, A => n1003, ZN => n999);
   U911 : AOI22_X1 port map( A1 => n940, A2 => n839, B1 => n1657, B2 => n381, 
                           ZN => n1003);
   U912 : NOR2_X1 port map( A1 => n1658, A2 => n1693, ZN => n940);
   U913 : AOI21_X1 port map( B1 => n1004, B2 => n1386, A => net74386, ZN => 
                           n997);
   U914 : AOI22_X1 port map( A1 => DATA1(12), A2 => net76217, B1 => net76297, 
                           B2 => n1756, ZN => n1004);
   U915 : OAI21_X1 port map( B1 => n1005, B2 => n1756, A => n1612_port, ZN => 
                           n996);
   U917 : NAND2_X1 port map( A1 => n1006, A2 => n1007, ZN => n995);
   U918 : AOI22_X1 port map( A1 => n1008, A2 => net82287, B1 => n1009, B2 => 
                           n350, ZN => n1007);
   U919 : OR2_X1 port map( A1 => n1010, A2 => n1011, ZN => n1009);
   U920 : OAI21_X1 port map( B1 => n1703, B2 => n1672, A => n1012, ZN => n1011)
                           ;
   U921 : AOI22_X1 port map( A1 => n357, A2 => n735, B1 => n356, B2 => n374, ZN
                           => n1012);
   U922 : OAI21_X1 port map( B1 => n1707, B2 => n1675, A => n1013, ZN => n1010)
                           ;
   U923 : AOI22_X1 port map( A1 => n519, A2 => n359, B1 => n456, B2 => n839, ZN
                           => n1013);
   U924 : OAI21_X1 port map( B1 => n1710, B2 => n1696, A => n1014, ZN => n1008)
                           ;
   U925 : AOI22_X1 port map( A1 => n1697, A2 => n1403, B1 => n576, B2 => n636, 
                           ZN => n1014);
   U926 : OAI21_X1 port map( B1 => n723, B2 => n1698, A => n1015, ZN => n485);
   U927 : NAND2_X1 port map( A1 => n1711, A2 => n1698, ZN => n1015);
   U928 : AOI22_X1 port map( A1 => N1622, A2 => net76325, B1 => N1991, B2 => 
                           n362, ZN => n1006);
   U930 : NAND2_X1 port map( A1 => net76617, A2 => n291, ZN => n1016);
   U933 : OAI21_X1 port map( B1 => n1432, B2 => n345, A => n1386, ZN => n1022);
   U934 : NAND2_X1 port map( A1 => n1023, A2 => n1024, ZN => n1021);
   U935 : OAI21_X1 port map( B1 => n1025, B2 => n1026, A => n1027, ZN => n1024)
                           ;
   U936 : OAI21_X1 port map( B1 => n684, B2 => n1658, A => n1028, ZN => n1026);
   U937 : AOI22_X1 port map( A1 => n1655, A2 => n438, B1 => n1656, B2 => n776, 
                           ZN => n1028);
   U938 : AOI21_X1 port map( B1 => n577, B2 => n1532, A => n1690, ZN => n684);
   U939 : AOI21_X1 port map( B1 => n1535, B2 => n774, A => n707, ZN => n1029);
   U940 : OAI21_X1 port map( B1 => net74284, B2 => net74295, A => n1030, ZN => 
                           n577);
   U941 : OAI21_X1 port map( B1 => n1721, B2 => n964, A => n1031, ZN => n1025);
   U942 : AOI21_X1 port map( B1 => n1652, B2 => n432, A => n418, ZN => n1031);
   U943 : AOI22_X1 port map( A1 => n397, A2 => n682, B1 => n1432, B2 => n1032, 
                           ZN => n1019);
   U944 : NAND2_X1 port map( A1 => n1033, A2 => net76311, ZN => n1032);
   U945 : AOI22_X1 port map( A1 => DATA1(10), A2 => net76217, B1 => net76297, 
                           B2 => net74264, ZN => n1033);
   U946 : NAND2_X1 port map( A1 => n1034, A2 => n1035, ZN => n682);
   U947 : AOI22_X1 port map( A1 => DATA1(9), A2 => n1582, B1 => DATA1(10), B2 
                           => n1561, ZN => n1035);
   U948 : AOI22_X1 port map( A1 => DATA1(7), A2 => n1573_port, B1 => DATA1(8), 
                           B2 => n1481, ZN => n1034);
   U949 : AOI22_X1 port map( A1 => n681, A2 => net82287, B1 => n1036, B2 => 
                           n350, ZN => n1018);
   U950 : OR2_X1 port map( A1 => n1037, A2 => n1038, ZN => n1036);
   U951 : OAI21_X1 port map( B1 => n1722, B2 => n1664, A => n1039, ZN => n1038)
                           ;
   U952 : AOI22_X1 port map( A1 => n356, A2 => n438, B1 => n357, B2 => n776, ZN
                           => n1039);
   U953 : NAND2_X1 port map( A1 => n1040, A2 => n1041, ZN => n776);
   U954 : AOI22_X1 port map( A1 => DATA1(22), A2 => n1582, B1 => DATA1(21), B2 
                           => n1475, ZN => n1041);
   U955 : AOI22_X1 port map( A1 => DATA1(24), A2 => n1573_port, B1 => DATA1(23)
                           , B2 => n1568_port, ZN => n1040);
   U956 : NAND2_X1 port map( A1 => n1042, A2 => n1043, ZN => n438);
   U957 : AOI22_X1 port map( A1 => DATA1(18), A2 => n1582, B1 => DATA1(17), B2 
                           => n1561, ZN => n1043);
   U958 : AOI22_X1 port map( A1 => DATA1(20), A2 => n1573_port, B1 => DATA1(19)
                           , B2 => n1481, ZN => n1042);
   U959 : NAND2_X1 port map( A1 => n1044, A2 => n1045, ZN => n774);
   U960 : AOI22_X1 port map( A1 => DATA1(26), A2 => n1582, B1 => DATA1(25), B2 
                           => n1475, ZN => n1045);
   U961 : AOI22_X1 port map( A1 => n1573_port, A2 => DATA1(28), B1 => DATA1(27)
                           , B2 => n1568_port, ZN => n1044);
   U962 : OAI21_X1 port map( B1 => n1721, B2 => n1672, A => n1046, ZN => n1037)
                           ;
   U963 : AOI22_X1 port map( A1 => n359, A2 => n578, B1 => n405, B2 => n432, ZN
                           => n1046);
   U964 : NAND2_X1 port map( A1 => n1047, A2 => n1048, ZN => n432);
   U965 : AOI22_X1 port map( A1 => DATA1(10), A2 => n1582, B1 => DATA1(9), B2 
                           => n1561, ZN => n1048);
   U966 : AOI22_X1 port map( A1 => DATA1(12), A2 => n1573_port, B1 => DATA1(11)
                           , B2 => n1481, ZN => n1047);
   U967 : OAI21_X1 port map( B1 => net74284, B2 => n1472, A => n1030, ZN => 
                           n578);
   U968 : AOI21_X1 port map( B1 => n1582, B2 => DATA1(30), A => n1049, ZN => 
                           n1030);
   U969 : NOR2_X1 port map( A1 => n1471, A2 => n1741, ZN => n1049);
   U970 : NAND2_X1 port map( A1 => n1050, A2 => n1051, ZN => n437);
   U971 : AOI22_X1 port map( A1 => DATA1(14), A2 => n1582, B1 => DATA1(13), B2 
                           => n1475, ZN => n1051);
   U972 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1573_port, B1 => DATA1(15)
                           , B2 => n1481, ZN => n1050);
   U973 : OAI21_X1 port map( B1 => n1701, B2 => n1696, A => n1052, ZN => n681);
   U974 : NAND2_X1 port map( A1 => n1540, A2 => n781, ZN => n1052);
   U975 : OAI21_X1 port map( B1 => n1472, B2 => n1767, A => n1053, ZN => n781);
   U976 : NOR2_X1 port map( A1 => n1054, A2 => n555, ZN => n1053);
   U977 : NOR2_X1 port map( A1 => n1765, A2 => n1471, ZN => n555);
   U978 : NAND2_X1 port map( A1 => n1055, A2 => n1056, ZN => n428);
   U979 : AOI21_X1 port map( B1 => DATA1(5), B2 => n518, A => n1057, ZN => 
                           n1056);
   U980 : AOI21_X1 port map( B1 => DATA1(6), B2 => n1475, A => n557, ZN => 
                           n1055);
   U981 : NOR2_X1 port map( A1 => n1763, A2 => n1472, ZN => n557);
   U982 : AOI22_X1 port map( A1 => N1620, A2 => net76325, B1 => N1989, B2 => 
                           n362, ZN => n1017);
   U983 : NOR4_X1 port map( A1 => n1058, A2 => n1059, A3 => n1060, A4 => n1061,
                           ZN => n292);
   U984 : AOI21_X1 port map( B1 => n1062, B2 => n1651, A => n1618_port, ZN => 
                           n1061);
   U985 : NOR2_X1 port map( A1 => n1620_port, A2 => net74248, ZN => n411);
   U986 : OAI21_X1 port map( B1 => n964, B2 => n1717, A => n1064, ZN => n1063);
   U987 : AOI21_X1 port map( B1 => n402, B2 => n1652, A => n418, ZN => n1064);
   U988 : NAND2_X1 port map( A1 => n1065, A2 => n1532, ZN => n964);
   U989 : AOI21_X1 port map( B1 => n445, B2 => n662, A => n1066, ZN => n1062);
   U990 : OAI21_X1 port map( B1 => n1719, B2 => n492, A => n1067, ZN => n1066);
   U991 : NAND2_X1 port map( A1 => n1656, A2 => n753, ZN => n1067);
   U992 : NAND2_X1 port map( A1 => n1065, A2 => n1538, ZN => n415);
   U993 : NAND2_X1 port map( A1 => n1065, A2 => n1540, ZN => n492);
   U994 : OAI21_X1 port map( B1 => n1068, B2 => n1696, A => n1069, ZN => n662);
   U995 : AOI21_X1 port map( B1 => n1535, B2 => n926, A => n707, ZN => n1069);
   U996 : NOR2_X1 port map( A1 => n1692, A2 => net74284, ZN => n707);
   U997 : NOR2_X1 port map( A1 => n1659, A2 => net74367, ZN => n445);
   U998 : AOI21_X1 port map( B1 => n1070, B2 => n1386, A => n1648, ZN => n1060)
                           ;
   U999 : AOI22_X1 port map( A1 => DATA1(11), A2 => net76217, B1 => net76297, 
                           B2 => n1757, ZN => n1070);
   U1000 : OAI21_X1 port map( B1 => n1720, B2 => n1668, A => n1071, ZN => n1059
                           );
   U1001 : AOI21_X1 port map( B1 => DATA1(11), B2 => n1072, A => n344, ZN => 
                           n1071);
   U1002 : NOR2_X1 port map( A1 => n1023, A2 => net74248, ZN => n344);
   U1003 : AOI21_X1 port map( B1 => n1073, B2 => DATA1(31), A => n1617_port, ZN
                           => n1023);
   U1004 : OAI21_X1 port map( B1 => n1450, B2 => n345, A => net76311, ZN => 
                           n1072);
   U1005 : NOR2_X1 port map( A1 => n1693, A2 => net74362, ZN => n397);
   U1006 : NAND2_X1 port map( A1 => n1074, A2 => n1075, ZN => n659);
   U1007 : AOI22_X1 port map( A1 => DATA1(10), A2 => n518, B1 => DATA1(11), B2 
                           => n1561, ZN => n1075);
   U1008 : AOI22_X1 port map( A1 => DATA1(8), A2 => n1573_port, B1 => DATA1(9),
                           B2 => n1481, ZN => n1074);
   U1009 : NAND2_X1 port map( A1 => n1076, A2 => n1077, ZN => n1058);
   U1010 : AOI22_X1 port map( A1 => n657, A2 => net82287, B1 => n1078, B2 => 
                           n350, ZN => n1077);
   U1011 : OR2_X1 port map( A1 => n1079, A2 => n1080, ZN => n1078);
   U1012 : OAI21_X1 port map( B1 => n1718, B2 => n1664, A => n1081, ZN => n1080
                           );
   U1013 : AOI22_X1 port map( A1 => n356, A2 => n409, B1 => n357, B2 => n753, 
                           ZN => n1081);
   U1014 : NAND2_X1 port map( A1 => n1082, A2 => n1083, ZN => n753);
   U1015 : AOI22_X1 port map( A1 => DATA1(23), A2 => n1582, B1 => DATA1(22), B2
                           => n1561, ZN => n1083);
   U1016 : AOI22_X1 port map( A1 => DATA1(25), A2 => n1573_port, B1 => 
                           DATA1(24), B2 => n1568_port, ZN => n1082);
   U1017 : NAND2_X1 port map( A1 => n1084, A2 => n1085, ZN => n409);
   U1018 : AOI22_X1 port map( A1 => DATA1(19), A2 => n1582, B1 => DATA1(18), B2
                           => n1561, ZN => n1085);
   U1019 : AOI22_X1 port map( A1 => DATA1(21), A2 => n1573_port, B1 => 
                           DATA1(20), B2 => n1481, ZN => n1084);
   U1020 : NAND2_X1 port map( A1 => n1086, A2 => n1087, ZN => n926);
   U1021 : AOI22_X1 port map( A1 => DATA1(27), A2 => n1582, B1 => DATA1(26), B2
                           => n1561, ZN => n1087);
   U1022 : AOI22_X1 port map( A1 => n1573_port, A2 => DATA1(29), B1 => 
                           n1568_port, B2 => DATA1(28), ZN => n1086);
   U1023 : OAI21_X1 port map( B1 => n1717, B2 => n1672, A => n1088, ZN => n1079
                           );
   U1024 : AOI22_X1 port map( A1 => n359, A2 => n1735, B1 => n405, B2 => n402, 
                           ZN => n1088);
   U1025 : NAND2_X1 port map( A1 => n1089, A2 => n1090, ZN => n402);
   U1026 : NOR2_X1 port map( A1 => n1091, A2 => n960, ZN => n1090);
   U1027 : NOR2_X1 port map( A1 => n1756, A2 => n1472, ZN => n960);
   U1028 : AOI22_X1 port map( A1 => DATA1(11), A2 => n1582, B1 => DATA1(10), B2
                           => n1475, ZN => n1089);
   U1029 : AOI21_X1 port map( B1 => DATA1(31), B2 => n1582, A => n591, ZN => 
                           n652);
   U1030 : NAND2_X1 port map( A1 => n1092, A2 => n1093, ZN => n408);
   U1031 : AOI22_X1 port map( A1 => DATA1(15), A2 => n1582, B1 => DATA1(14), B2
                           => n1475, ZN => n1093);
   U1032 : AOI22_X1 port map( A1 => DATA1(17), A2 => n1573_port, B1 => 
                           DATA1(16), B2 => n1481, ZN => n1092);
   U1034 : OAI21_X1 port map( B1 => n1716, B2 => n1688, A => n1096, ZN => n657)
                           ;
   U1035 : NAND2_X1 port map( A1 => n1532, A2 => n398, ZN => n1096);
   U1036 : NAND2_X1 port map( A1 => n1097, A2 => n1098, ZN => n398);
   U1037 : AOI22_X1 port map( A1 => DATA1(6), A2 => n1582, B1 => DATA1(7), B2 
                           => n1561, ZN => n1098);
   U1038 : AOI22_X1 port map( A1 => DATA1(4), A2 => n1573_port, B1 => DATA1(5),
                           B2 => n1481, ZN => n1097);
   U1039 : NAND2_X1 port map( A1 => n1099, A2 => n1100, ZN => n566);
   U1040 : AOI22_X1 port map( A1 => n1461, A2 => n1582, B1 => n1404, B2 => 
                           n1561, ZN => n1100);
   U1041 : AOI22_X1 port map( A1 => n1399, A2 => n1573_port, B1 => n1405, B2 =>
                           n1481, ZN => n1099);
   U1042 : AOI22_X1 port map( A1 => N1621, A2 => net76325, B1 => N1990, B2 => 
                           n362, ZN => n1076);
   U1043 : OAI21_X1 port map( B1 => n289, B2 => net76321, A => n1101, ZN => 
                           OUTALU(0));
   U1044 : NAND2_X1 port map( A1 => n268, A2 => net74246, ZN => n1101);
   U1045 : NAND2_X1 port map( A1 => n1102, A2 => n1103, ZN => n268);
   U1046 : NOR4_X1 port map( A1 => n544, A2 => n1104, A3 => n1105, A4 => n1106,
                           ZN => n1103);
   U1047 : AOI21_X1 port map( B1 => n1107, B2 => n1386, A => net74295, ZN => 
                           n1106);
   U1048 : AOI22_X1 port map( A1 => n1405, A2 => n341, B1 => n1385, B2 => n1766
                           , ZN => n1107);
   U1049 : OAI21_X1 port map( B1 => net82639, B2 => n1108, A => n1109, ZN => 
                           n341);
   U1050 : NOR2_X1 port map( A1 => n1110, A2 => n1766, ZN => n1105);
   U1052 : OAI21_X1 port map( B1 => net74243, B2 => n1094, A => n1111, ZN => 
                           n488);
   U1053 : OR2_X1 port map( A1 => n1109, A2 => net92255, ZN => n1111);
   U1054 : NAND2_X1 port map( A1 => n301, A2 => n1112, ZN => n1109);
   U1055 : NAND2_X1 port map( A1 => n301, A2 => n1113, ZN => n345);
   U1056 : OAI21_X1 port map( B1 => net76624, B2 => n1114, A => net74236, ZN =>
                           n1113);
   U1057 : AOI21_X1 port map( B1 => net74247, B2 => n546, A => n1115, ZN => 
                           n1104);
   U1058 : NOR4_X1 port map( A1 => n1116, A2 => n1661, A3 => n1117, A4 => n1118
                           , ZN => n1115);
   U1059 : NOR2_X1 port map( A1 => n1119, A2 => n1675, ZN => n1118);
   U1060 : NOR4_X1 port map( A1 => n1054, A2 => n723, A3 => n1057, A4 => n1120,
                           ZN => n1119);
   U1061 : NOR2_X1 port map( A1 => n1472, A2 => n1765, ZN => n1120);
   U1062 : NOR2_X1 port map( A1 => n1764, A2 => n1577_port, ZN => n1057);
   U1063 : NOR2_X1 port map( A1 => n1766, A2 => n1585, ZN => n1054);
   U1064 : NOR2_X1 port map( A1 => n885, A2 => net74367, ZN => n1117);
   U1065 : AOI21_X1 port map( B1 => n360, B2 => n1538, A => n1121, ZN => n885);
   U1066 : NOR2_X1 port map( A1 => n1688, A2 => n1715, ZN => n1121);
   U1067 : NAND2_X1 port map( A1 => n1122, A2 => n1123, ZN => n460);
   U1068 : AOI22_X1 port map( A1 => DATA1(25), A2 => n1582, B1 => DATA1(24), B2
                           => n1475, ZN => n1123);
   U1069 : AOI22_X1 port map( A1 => DATA1(27), A2 => n1573_port, B1 => 
                           DATA1(26), B2 => n1568_port, ZN => n1122);
   U1070 : NAND2_X1 port map( A1 => n1124, A2 => n1125, ZN => n360);
   U1071 : AOI22_X1 port map( A1 => DATA1(29), A2 => n1582, B1 => DATA1(28), B2
                           => n1475, ZN => n1125);
   U1072 : AOI22_X1 port map( A1 => n1573_port, A2 => DATA1(31), B1 => 
                           DATA1(30), B2 => n1568_port, ZN => n1124);
   U1073 : AOI21_X1 port map( B1 => n337, B2 => n1545, A => n1127, ZN => n1126)
                           ;
   U1074 : NOR2_X1 port map( A1 => n1662, A2 => n1700, ZN => n1127);
   U1075 : NAND2_X1 port map( A1 => n1128, A2 => n1129, ZN => n336);
   U1076 : AOI22_X1 port map( A1 => DATA1(21), A2 => n1582, B1 => DATA1(20), B2
                           => n1561, ZN => n1129);
   U1077 : NOR2_X1 port map( A1 => n691, A2 => n1130, ZN => n1128);
   U1078 : NOR2_X1 port map( A1 => n1746, A2 => n1577_port, ZN => n691);
   U1079 : NAND2_X1 port map( A1 => n1131, A2 => n1132, ZN => n337);
   U1080 : AOI22_X1 port map( A1 => DATA1(13), A2 => n1582, B1 => DATA1(12), B2
                           => n1561, ZN => n1132);
   U1081 : AOI22_X1 port map( A1 => DATA1(15), A2 => n1573_port, B1 => 
                           DATA1(14), B2 => n1481, ZN => n1131);
   U1082 : OAI21_X1 port map( B1 => n1713, B2 => n1669, A => n1133, ZN => n1116
                           );
   U1083 : AOI22_X1 port map( A1 => n361, A2 => n461, B1 => n456, B2 => n335, 
                           ZN => n1133);
   U1084 : NAND2_X1 port map( A1 => n1134, A2 => n1135, ZN => n335);
   U1085 : AOI22_X1 port map( A1 => DATA1(17), A2 => n1582, B1 => DATA1(16), B2
                           => n1561, ZN => n1135);
   U1086 : AOI22_X1 port map( A1 => DATA1(19), A2 => n1573_port, B1 => 
                           DATA1(18), B2 => n1481, ZN => n1134);
   U1087 : NAND2_X1 port map( A1 => n1136, A2 => n1137, ZN => n461);
   U1088 : AOI21_X1 port map( B1 => DATA1(5), B2 => n1582, A => n1138, ZN => 
                           n1137);
   U1089 : AOI22_X1 port map( A1 => DATA1(7), A2 => n1573_port, B1 => DATA1(6),
                           B2 => n1568_port, ZN => n1136);
   U1090 : NAND2_X1 port map( A1 => n1139, A2 => n1140, ZN => n473);
   U1091 : AOI22_X1 port map( A1 => DATA1(9), A2 => n1582, B1 => DATA1(8), B2 
                           => n1561, ZN => n1140);
   U1092 : AOI22_X1 port map( A1 => DATA1(11), A2 => n1573_port, B1 => 
                           DATA1(10), B2 => n1568_port, ZN => n1139);
   U1093 : NAND2_X1 port map( A1 => n1141, A2 => n1142, ZN => n546);
   U1094 : NOR2_X1 port map( A1 => net74248, A2 => n1779, ZN => n1141);
   U1096 : NAND2_X1 port map( A1 => n1144, A2 => n315, ZN => n1143);
   U1098 : NOR2_X1 port map( A1 => net74248, A2 => n1146, ZN => n544);
   U1099 : NOR4_X1 port map( A1 => n1625_port, A2 => n1147, A3 => n1148, A4 => 
                           n1149, ZN => n1146);
   U1100 : AOI21_X1 port map( B1 => N1980, B2 => n362, A => n1150, ZN => n1102)
                           ;
   U1101 : OAI21_X1 port map( B1 => n462, B2 => n1673, A => n1151, ZN => n1150)
                           ;
   U1102 : NAND2_X1 port map( A1 => N1611, A2 => net76327, ZN => n1151);
   U1103 : NOR2_X1 port map( A1 => n1675, A2 => net74250, ZN => n514);
   U1104 : NOR2_X1 port map( A1 => n1152, A2 => n818, ZN => n462);
   U1105 : NOR2_X1 port map( A1 => n1766, A2 => n1471, ZN => n818);
   U1108 : AOI21_X1 port map( B1 => n1155, B2 => n1156, A => n1157, ZN => n1154
                           );
   U1110 : NOR3_X1 port map( A1 => n528, A2 => n302, A3 => n1159, ZN => n1153);
   U1111 : OAI21_X1 port map( B1 => n1161, B2 => n1160, A => n1162, ZN => NEG);
   U1112 : NAND2_X1 port map( A1 => n1157, A2 => N2010, ZN => n1162);
   U1113 : OAI33_X1 port map( A1 => n1163, A2 => n1357, A3 => net74231, B1 => 
                           n1164, B2 => net82773, B3 => net74455, ZN => n1161);
   U1115 : NOR2_X1 port map( A1 => n311, A2 => n1770, ZN => n1165);
   U1117 : OAI21_X1 port map( B1 => n1168, B2 => n1169, A => n1170, ZN => n1167
                           );
   U1119 : NOR2_X1 port map( A1 => net74235, A2 => net88905, ZN => n1169);
   U1121 : NAND2_X1 port map( A1 => n302, A2 => net83941, ZN => n1166);
   U1123 : OAI21_X1 port map( B1 => net83085, B2 => n1373, A => n1173, ZN => 
                           n1163);
   U1127 : OAI21_X1 port map( B1 => n576, B2 => net74284, A => n909, ZN => 
                           n1176);
   U1128 : NOR4_X1 port map( A1 => n1617_port, A2 => n1147, A3 => n1177, A4 => 
                           n1148, ZN => n909);
   U1129 : OAI21_X1 port map( B1 => net74284, B2 => n1638_port, A => n1178, ZN 
                           => n1148);
   U1130 : AOI21_X1 port map( B1 => n1179, B2 => net74367, A => net74284, ZN =>
                           n1177);
   U1131 : OAI21_X1 port map( B1 => n1641_port, B2 => net74284, A => n1660, ZN 
                           => n1147);
   U1132 : NOR2_X1 port map( A1 => net74284, A2 => n1180, ZN => n418);
   U1133 : NAND2_X1 port map( A1 => n1535, A2 => n1734, ZN => n1175);
   U1134 : AOI21_X1 port map( B1 => n1471, B2 => DATA1(31), A => n591, ZN => 
                           n1068);
   U1135 : NOR2_X1 port map( A1 => n1740, A2 => n1471, ZN => n591);
   U1136 : NAND2_X1 port map( A1 => n1183, A2 => n1065, ZN => n904);
   U1137 : NOR2_X1 port map( A1 => n1181, A2 => n1779, ZN => n1183);
   U1139 : AOI21_X1 port map( B1 => n1187, B2 => n1155, A => n1188, ZN => n1160
                           );
   U1141 : NAND2_X1 port map( A1 => net76624, A2 => net83091, ZN => n1189);
   U1142 : AOI21_X1 port map( B1 => n1190, B2 => n1191, A => n1769, ZN => n1187
                           );
   U1143 : OAI21_X1 port map( B1 => net74238, B2 => net83941, A => net86253, ZN
                           => n1190);
   U1145 : NAND2_X1 port map( A1 => n1467, A2 => net76617, ZN => n1193);
   U1148 : AOI21_X1 port map( B1 => n1155, B2 => n1201, A => n1157, ZN => n1200
                           );
   U1152 : OAI21_X1 port map( B1 => net76624, B2 => net74229, A => n1158, ZN =>
                           n1201);
   U1155 : NOR2_X1 port map( A1 => net74238, A2 => net74226, ZN => n302);
   U1156 : OR2_X1 port map( A1 => n528, A2 => n1159, ZN => n1204);
   U1157 : NOR2_X1 port map( A1 => n1205, A2 => net74238, ZN => n1159);
   U1158 : OR2_X1 port map( A1 => net82733, A2 => n311, ZN => n1205);
   U1159 : NAND2_X1 port map( A1 => n1206, A2 => n313, ZN => n528);
   U1161 : AOI22_X1 port map( A1 => n1145, A2 => net92271, B1 => n315, B2 => 
                           n1208, ZN => n1207);
   U1162 : NOR2_X1 port map( A1 => n1471, A2 => net74284, ZN => n519);
   U1164 : NAND2_X1 port map( A1 => n1209, A2 => n301, ZN => n510);
   U1165 : NOR2_X1 port map( A1 => net77046, A2 => net83926, ZN => n301);
   U1166 : NOR2_X1 port map( A1 => net92255, A2 => n1114, ZN => n1209);
   U1167 : OAI21_X1 port map( B1 => net74248, B2 => net74284, A => n1210, ZN =>
                           n1195);
   U1168 : OAI21_X1 port map( B1 => n1211, B2 => n1212, A => n582, ZN => n1210)
                           ;
   U1170 : OR2_X1 port map( A1 => n1094, A2 => net82639, ZN => n1213);
   U1171 : NAND2_X1 port map( A1 => n1214, A2 => n1112, ZN => n1095);
   U1172 : NOR2_X1 port map( A1 => n1191, A2 => net82733, ZN => n1112);
   U1173 : NOR2_X1 port map( A1 => net83085, A2 => net76624, ZN => n1214);
   U1174 : OAI21_X1 port map( B1 => n1712, B2 => n1669, A => n1215, ZN => n1212
                           );
   U1175 : AOI22_X1 port map( A1 => n357, A2 => n642, B1 => n456, B2 => n635, 
                           ZN => n1215);
   U1176 : NAND2_X1 port map( A1 => n1216, A2 => n1217, ZN => n635);
   U1177 : AOI21_X1 port map( B1 => DATA1(15), B2 => n1582, A => n1091, ZN => 
                           n1217);
   U1178 : NOR2_X1 port map( A1 => n1755, A2 => n1577_port, ZN => n1091);
   U1179 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1475, B1 => DATA1(14), B2
                           => n1481, ZN => n1216);
   U1180 : NAND2_X1 port map( A1 => n1218, A2 => n1219, ZN => n642);
   U1181 : AOI22_X1 port map( A1 => DATA1(19), A2 => n1582, B1 => DATA1(20), B2
                           => n1561, ZN => n1219);
   U1182 : AOI22_X1 port map( A1 => DATA1(17), A2 => n1573_port, B1 => 
                           DATA1(18), B2 => n1568_port, ZN => n1218);
   U1183 : NAND2_X1 port map( A1 => n1220, A2 => n1221, ZN => n733);
   U1184 : AOI21_X1 port map( B1 => DATA1(23), B2 => n1582, A => n1130, ZN => 
                           n1221);
   U1185 : NOR2_X1 port map( A1 => n1747, A2 => n1472, ZN => n1130);
   U1186 : AOI22_X1 port map( A1 => DATA1(24), A2 => n1561, B1 => DATA1(21), B2
                           => n1573_port, ZN => n1220);
   U1187 : NAND2_X1 port map( A1 => n1222, A2 => n1223, ZN => n1211);
   U1188 : AOI22_X1 port map( A1 => net76732, A2 => n1224, B1 => n405, B2 => 
                           n1225, ZN => n1223);
   U1189 : OAI21_X1 port map( B1 => n1472, B2 => n1740, A => n1226, ZN => n1225
                           );
   U1190 : AOI22_X1 port map( A1 => n1582, A2 => DATA1(31), B1 => n1573_port, 
                           B2 => DATA1(29), ZN => n1226);
   U1191 : OAI21_X1 port map( B1 => n1710, B2 => n1688, A => n1227, ZN => n1224
                           );
   U1192 : NAND2_X1 port map( A1 => n1538, A2 => n725, ZN => n1227);
   U1193 : NAND2_X1 port map( A1 => n1228, A2 => n1229, ZN => n725);
   U1194 : AOI21_X1 port map( B1 => n1405, B2 => n1573_port, A => n1138, ZN => 
                           n1229);
   U1195 : NOR2_X1 port map( A1 => n1763, A2 => n1471, ZN => n1138);
   U1196 : AOI21_X1 port map( B1 => n1461, B2 => n1481, A => n556, ZN => n1228)
                           ;
   U1197 : NOR2_X1 port map( A1 => n1764, A2 => n1585, ZN => n556);
   U1198 : NAND2_X1 port map( A1 => n1230, A2 => n1231, ZN => n639);
   U1199 : AOI22_X1 port map( A1 => DATA1(7), A2 => n518, B1 => DATA1(8), B2 =>
                           n1561, ZN => n1231);
   U1200 : AOI22_X1 port map( A1 => DATA1(5), A2 => n1573_port, B1 => DATA1(6),
                           B2 => n1568_port, ZN => n1230);
   U1201 : AOI22_X1 port map( A1 => n359, A2 => n636, B1 => n361, B2 => n641, 
                           ZN => n1222);
   U1202 : NAND2_X1 port map( A1 => n1232, A2 => n1233, ZN => n641);
   U1203 : AOI22_X1 port map( A1 => DATA1(27), A2 => n1582, B1 => DATA1(28), B2
                           => n1561, ZN => n1233);
   U1204 : AOI22_X1 port map( A1 => DATA1(25), A2 => n1573_port, B1 => 
                           DATA1(26), B2 => n1568_port, ZN => n1232);
   U1205 : NAND2_X1 port map( A1 => n1234, A2 => n1235, ZN => n636);
   U1206 : AOI22_X1 port map( A1 => DATA1(11), A2 => n1582, B1 => DATA1(12), B2
                           => n1561, ZN => n1235);
   U1207 : AOI22_X1 port map( A1 => DATA1(9), A2 => n1573_port, B1 => DATA1(10)
                           , B2 => n1568_port, ZN => n1234);
   U1211 : NOR2_X1 port map( A1 => n1239, A2 => n1240, ZN => n289);
   U1212 : OAI21_X1 port map( B1 => n1241, B2 => net82639, A => n1242, ZN => 
                           n1240);
   U1213 : AOI22_X1 port map( A1 => n1155, A2 => n1243, B1 => N1610, B2 => 
                           net76327, ZN => n1242);
   U1216 : OR2_X1 port map( A1 => n1245, A2 => n1246, ZN => n1243);
   U1217 : OAI21_X1 port map( B1 => N1577, B2 => n1094, A => n1247, ZN => n1246
                           );
   U1218 : AOI22_X1 port map( A1 => N1576, A2 => net74234, B1 => n1145, B2 => 
                           net74464, ZN => n1247);
   U1219 : OAI21_X1 port map( B1 => net74463, B2 => n313, A => n1248, ZN => 
                           n1245);
   U1220 : AOI21_X1 port map( B1 => N1979, B2 => n1249, A => n1250, ZN => n1248
                           );
   U1221 : NOR3_X1 port map( A1 => net74225, A2 => n1588, A3 => net74238, ZN =>
                           n1250);
   U1223 : OAI21_X1 port map( B1 => net92259, B2 => n251, A => n1192, ZN => 
                           n1158);
   U1224 : NAND2_X1 port map( A1 => n1253, A2 => net92259, ZN => n1192);
   U1226 : NAND2_X1 port map( A1 => net92259, A2 => n320, ZN => n1252);
   U1228 : NOR3_X1 port map( A1 => n1254, A2 => n1255, A3 => n1256, ZN => n1241
                           );
   U1229 : OAI33_X1 port map( A1 => n1733, A2 => n1675, A3 => n1094, B1 => 
                           n1108, B2 => n1738, B3 => n1767, ZN => n1256);
   U1230 : NAND2_X1 port map( A1 => n251, A2 => net92254, ZN => n1108);
   U1231 : NAND2_X1 port map( A1 => n1257, A2 => n310, ZN => n1094);
   U1232 : AOI21_X1 port map( B1 => n1206, B2 => n313, A => n1737, ZN => n1255)
                           ;
   U1233 : NAND2_X1 port map( A1 => n314, A2 => net92254, ZN => n313);
   U1234 : OAI21_X1 port map( B1 => n1258, B2 => n1236, A => n1259, ZN => n1254
                           );
   U1235 : NAND2_X1 port map( A1 => n1145, A2 => n1260, ZN => n1259);
   U1236 : NOR2_X1 port map( A1 => net74225, A2 => net74235, ZN => n1145);
   U1238 : NAND2_X1 port map( A1 => n1257, A2 => n314, ZN => n1236);
   U1239 : NOR2_X1 port map( A1 => net92259, A2 => net76624, ZN => n1257);
   U1240 : OAI21_X1 port map( B1 => n1261, B2 => net74238, A => n1262, ZN => 
                           n1239);
   U1244 : OAI21_X1 port map( B1 => n1266, B2 => n1267, A => ALU_OPCODE(0), ZN 
                           => n1265);
   U1245 : NOR2_X1 port map( A1 => n1268, A2 => net77046, ZN => n1267);
   U1246 : AOI21_X1 port map( B1 => n321, B2 => net74464, A => n1269, ZN => 
                           n1268);
   U1248 : NOR3_X1 port map( A1 => n1270, A2 => net83085, A3 => n321, ZN => 
                           n1266);
   U1249 : NOR2_X1 port map( A1 => net82733, A2 => net76624, ZN => n321);
   U1250 : AOI22_X1 port map( A1 => N1979, A2 => net74226, B1 => net86253, B2 
                           => net74463, ZN => n1270);
   U1252 : AOI21_X1 port map( B1 => n1271, B2 => n1272, A => net83926, ZN => 
                           n1263);
   U1254 : OAI21_X1 port map( B1 => net76624, B2 => n1275, A => n1276, ZN => 
                           n1273);
   U1255 : AOI22_X1 port map( A1 => n251, A2 => n1251, B1 => n314, B2 => n1277,
                           ZN => n1271);
   U1256 : OAI21_X1 port map( B1 => net76624, B2 => n1589, A => n1278, ZN => 
                           n1251);
   U1257 : NAND2_X1 port map( A1 => N1573, A2 => net76624, ZN => n1278);
   U1258 : AOI21_X1 port map( B1 => n1279, B2 => n315, A => n1280, ZN => n1261)
                           ;
   U1259 : AOI21_X1 port map( B1 => n1281, B2 => n1282, A => net83926, ZN => 
                           n1280);
   U1260 : OAI21_X1 port map( B1 => n1283, B2 => n251, A => N1979, ZN => n1282)
                           ;
   U1261 : NOR3_X1 port map( A1 => n311, A2 => net83085, A3 => net82733, ZN => 
                           n1283);
   U1262 : XNOR2_X1 port map( A => net76624, B => n1284, ZN => n311);
   U1263 : NOR4_X1 port map( A1 => DATA2(31), A2 => n1471, A3 => n333, A4 => 
                           n1620_port, ZN => n1284);
   U1264 : NOR2_X1 port map( A1 => n1073, A2 => n1185, ZN => n1027);
   U1266 : NOR3_X1 port map( A1 => DATA2(19), A2 => DATA2(21), A3 => DATA2(20),
                           ZN => n1288);
   U1267 : NOR3_X1 port map( A1 => n1448, A2 => DATA2(18), A3 => n1438, ZN => 
                           n1287);
   U1268 : NOR3_X1 port map( A1 => n1629_port, A2 => n1450, A3 => net83048, ZN 
                           => n1286);
   U1269 : NOR3_X1 port map( A1 => n1624_port, A2 => n1290, A3 => n1291, ZN => 
                           n1285);
   U1270 : NOR4_X1 port map( A1 => DATA2(28), A2 => DATA2(27), A3 => DATA2(26),
                           A4 => DATA2(25), ZN => n1179);
   U1271 : NAND2_X1 port map( A1 => n1065, A2 => n1535, ZN => n333);
   U1272 : NOR2_X1 port map( A1 => n1659, A2 => net76732, ZN => n1065);
   U1273 : OAI21_X1 port map( B1 => n1292, B2 => n1293, A => net83085, ZN => 
                           n1281);
   U1274 : NOR2_X1 port map( A1 => n1294, A2 => net74225, ZN => n1293);
   U1275 : AOI22_X1 port map( A1 => net76624, A2 => n1739, B1 => n1399, B2 => 
                           DATA2(0), ZN => n1294);
   U1276 : NOR2_X1 port map( A1 => DATA2(0), A2 => n1399, ZN => n1275);
   U1277 : NOR3_X1 port map( A1 => net74224, A2 => net76624, A3 => n1276, ZN =>
                           n1292);
   U1278 : XNOR2_X1 port map( A => n1399, B => DATA2(0), ZN => n1276);
   U1280 : AOI21_X1 port map( B1 => n1295, B2 => n1296, A => net83085, ZN => 
                           n1279);
   U1281 : AOI21_X1 port map( B1 => n1297, B2 => n314, A => n1298, ZN => n1296)
                           ;
   U1282 : NOR2_X1 port map( A1 => net76624, A2 => n1299, ZN => n1298);
   U1283 : AOI21_X1 port map( B1 => n314, B2 => n1260, A => n1300, ZN => n1299)
                           ;
   U1284 : NOR3_X1 port map( A1 => n1733, A2 => n1675, A3 => net74225, ZN => 
                           n1300);
   U1285 : NOR2_X1 port map( A1 => net86253, A2 => net82733, ZN => n310);
   U1286 : NOR2_X1 port map( A1 => n1767, A2 => n1471, ZN => n723);
   U1288 : NOR2_X1 port map( A1 => n1258, A2 => net83941, ZN => n1297);
   U1289 : NOR2_X1 port map( A1 => n1301, A2 => n1149, ZN => n1258);
   U1290 : NAND2_X1 port map( A1 => n1302, A2 => n1182, ZN => n1149);
   U1291 : NAND2_X1 port map( A1 => DATA1(31), A2 => n1185, ZN => n1182);
   U1292 : OAI21_X1 port map( B1 => DATA2(28), B2 => DATA2(27), A => DATA1(31),
                           ZN => n1302);
   U1293 : NOR4_X1 port map( A1 => DATA2(28), A2 => DATA2(27), A3 => n1303, A4 
                           => n1185, ZN => n1301);
   U1294 : OR2_X1 port map( A1 => DATA2(29), A2 => DATA2(30), ZN => n1185);
   U1295 : NOR3_X1 port map( A1 => n1625_port, A2 => n1630_port, A3 => n1304, 
                           ZN => n1303);
   U1296 : NOR4_X1 port map( A1 => DATA2(26), A2 => DATA2(25), A3 => n1305, A4 
                           => n1186, ZN => n1304);
   U1297 : AOI22_X1 port map( A1 => DATA1(31), A2 => n1306, B1 => n1637_port, 
                           B2 => n1260, ZN => n1305);
   U1298 : OR2_X1 port map( A1 => n1307, A2 => n1308, ZN => n1260);
   U1299 : OAI21_X1 port map( B1 => n1706, B2 => n1672, A => n1309, ZN => n1308
                           );
   U1300 : AOI22_X1 port map( A1 => n1545, A2 => n491, B1 => n1549, B2 => n376,
                           ZN => n1309);
   U1301 : NAND2_X1 port map( A1 => n1310, A2 => n1311, ZN => n376);
   U1302 : AOI22_X1 port map( A1 => DATA1(8), A2 => n518, B1 => DATA1(7), B2 =>
                           n1561, ZN => n1311);
   U1303 : AOI22_X1 port map( A1 => DATA1(10), A2 => n520, B1 => DATA1(9), B2 
                           => n1568_port, ZN => n1310);
   U1304 : NOR2_X1 port map( A1 => n1688, A2 => net76732, ZN => n356);
   U1305 : NAND2_X1 port map( A1 => n1312, A2 => n1313, ZN => n491);
   U1306 : AOI22_X1 port map( A1 => DATA1(12), A2 => n518, B1 => DATA1(11), B2 
                           => n1561, ZN => n1313);
   U1307 : AOI22_X1 port map( A1 => DATA1(14), A2 => n520, B1 => DATA1(13), B2 
                           => n1568_port, ZN => n1312);
   U1308 : NOR2_X1 port map( A1 => n1679, A2 => net76732, ZN => n357);
   U1309 : NOR2_X1 port map( A1 => n1696, A2 => net76732, ZN => n361);
   U1310 : NAND2_X1 port map( A1 => n1314, A2 => n1315, ZN => n498);
   U1311 : AOI22_X1 port map( A1 => DATA1(4), A2 => n518, B1 => n1404, B2 => 
                           n1561, ZN => n1315);
   U1312 : AOI22_X1 port map( A1 => DATA1(6), A2 => n520, B1 => DATA1(5), B2 =>
                           n1568_port, ZN => n1314);
   U1313 : NAND2_X1 port map( A1 => n1316, A2 => n1317, ZN => n1307);
   U1314 : AOI22_X1 port map( A1 => net76732, A2 => n905, B1 => n405, B2 => 
                           n1318, ZN => n1317);
   U1315 : OAI21_X1 port map( B1 => n1472, B2 => n1766, A => n1319, ZN => n1318
                           );
   U1316 : AOI21_X1 port map( B1 => n1461, B2 => n520, A => n1152, ZN => n1319)
                           ;
   U1317 : NOR2_X1 port map( A1 => n1767, A2 => n1585, ZN => n1152);
   U1318 : NOR2_X1 port map( A1 => n1693, A2 => net76732, ZN => n405);
   U1319 : OAI21_X1 port map( B1 => n1704, B2 => n1679, A => n1320, ZN => n905)
                           ;
   U1320 : NAND2_X1 port map( A1 => n1540, A2 => n735, ZN => n1320);
   U1321 : NAND2_X1 port map( A1 => n1321, A2 => n1322, ZN => n735);
   U1322 : AOI22_X1 port map( A1 => DATA1(24), A2 => n518, B1 => DATA1(23), B2 
                           => n1561, ZN => n1322);
   U1323 : AOI22_X1 port map( A1 => DATA1(26), A2 => n520, B1 => DATA1(25), B2 
                           => n1568_port, ZN => n1321);
   U1324 : NOR2_X1 port map( A1 => n1692, A2 => DATA2(2), ZN => n562);
   U1325 : NOR2_X1 port map( A1 => n1692, A2 => n1698, ZN => n563);
   U1326 : NAND2_X1 port map( A1 => n1323, A2 => n1324, ZN => n839);
   U1327 : AOI22_X1 port map( A1 => DATA1(28), A2 => n518, B1 => DATA1(27), B2 
                           => n1561, ZN => n1324);
   U1328 : AOI22_X1 port map( A1 => DATA1(30), A2 => n520, B1 => n1568_port, B2
                           => DATA1(29), ZN => n1323);
   U1329 : AOI22_X1 port map( A1 => n359, A2 => n374, B1 => n456, B2 => n381, 
                           ZN => n1316);
   U1330 : NAND2_X1 port map( A1 => n1325, A2 => n1326, ZN => n381);
   U1331 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1582, B1 => DATA1(15), B2
                           => n1561, ZN => n1326);
   U1332 : AOI22_X1 port map( A1 => DATA1(18), A2 => n520, B1 => DATA1(17), B2 
                           => n1568_port, ZN => n1325);
   U1333 : NOR2_X1 port map( A1 => n1693, A2 => net74367, ZN => n456);
   U1334 : NOR2_X1 port map( A1 => n1403, A2 => DATA2(2), ZN => n576);
   U1335 : NAND2_X1 port map( A1 => n1327, A2 => n1328, ZN => n374);
   U1336 : AOI22_X1 port map( A1 => DATA1(20), A2 => n1582, B1 => DATA1(19), B2
                           => n1561, ZN => n1328);
   U1338 : NOR2_X1 port map( A1 => n1738, A2 => DATA2(1), ZN => n518);
   U1339 : AOI22_X1 port map( A1 => DATA1(22), A2 => n520, B1 => DATA1(21), B2 
                           => n1568_port, ZN => n1327);
   U1341 : NOR2_X1 port map( A1 => net74295, A2 => n1738, ZN => n520);
   U1342 : NOR2_X1 port map( A1 => n1696, A2 => net74367, ZN => n359);
   U1343 : NOR2_X1 port map( A1 => n1698, A2 => n1403, ZN => n465);
   U1344 : NAND2_X1 port map( A1 => n1142, A2 => n1638_port, ZN => n1306);
   U1345 : NOR2_X1 port map( A1 => n1659, A2 => n1181, ZN => n1142);
   U1346 : NAND2_X1 port map( A1 => n1329, A2 => n1330, ZN => n1181);
   U1347 : NOR4_X1 port map( A1 => DATA2(18), A2 => n1438, A3 => n1448, A4 => 
                           net83048, ZN => n1330);
   U1348 : NOR3_X1 port map( A1 => n1291, A2 => n1450, A3 => n1290, ZN => n1329
                           );
   U1349 : NAND2_X1 port map( A1 => n1331, A2 => n1646, ZN => n1290);
   U1350 : NOR2_X1 port map( A1 => DATA2(17), A2 => DATA2(16), ZN => n1331);
   U1351 : NAND2_X1 port map( A1 => n1332, A2 => n1649, ZN => n1291);
   U1352 : NOR2_X1 port map( A1 => n1416, A2 => n1460, ZN => n1332);
   U1353 : NOR2_X1 port map( A1 => n1333, A2 => n1456, ZN => n1180);
   U1354 : OR2_X1 port map( A1 => n1457, A2 => net82473, ZN => n1333);
   U1355 : NAND2_X1 port map( A1 => DATA1(31), A2 => n1186, ZN => n1178);
   U1356 : NAND2_X1 port map( A1 => n1334, A2 => n1289, ZN => n1186);
   U1357 : NOR2_X1 port map( A1 => n1335, A2 => DATA2(22), ZN => n1289);
   U1358 : OR2_X1 port map( A1 => DATA2(24), A2 => DATA2(23), ZN => n1335);
   U1359 : NOR2_X1 port map( A1 => DATA2(21), A2 => DATA2(20), ZN => n1334);
   U1360 : OAI21_X1 port map( B1 => DATA2(26), B2 => DATA2(25), A => DATA1(31),
                           ZN => n1336);
   U1362 : XNOR2_X1 port map( A => net83941, B => N1568, ZN => n1277);
   U1365 : AOI21_X1 port map( B1 => net83941, B2 => N1573, A => n1337, ZN => 
                           n1274);
   U1366 : NOR2_X1 port map( A1 => n1589, A2 => net83941, ZN => n1337);
   U1126 : OAI21_X1 port map( B1 => n904, B2 => n1175, A => net74426, ZN => 
                           n509);
   U1140 : OAI21_X1 port map( B1 => net74233, B2 => n1189, A => net82639, ZN =>
                           n1188);
   U1097 : NOR2_X1 port map( A1 => net76624, A2 => net74233, ZN => n1144);
   U279 : AOI22_X1 port map( A1 => n305, A2 => net74231, B1 => n306, B2 => n307
                           , ZN => n304);
   U1372 : NOR2_X1 port map( A1 => n1114, A2 => net83085, ZN => n1208);
   U1373 : OR2_X1 port map( A1 => n1191, A2 => net82508, ZN => n1114);
   U255 : NAND2_X1 port map( A1 => n251, A2 => net92255, ZN => n250);
   U1125 : AOI21_X1 port map( B1 => net74238, B2 => net82508, A => net77046, ZN
                           => n1174);
   U1222 : OAI21_X1 port map( B1 => net82508, B2 => n1252, A => n1158, ZN => 
                           n1249);
   U1247 : OAI33_X1 port map( A1 => net74464, A2 => net82733, A3 => net83941, 
                           B1 => net74463, B2 => net76624, B3 => net82508, ZN 
                           => n1269);
   U1371 : XNOR2_X1 port map( A => net82733, B => net92255, ZN => n320);
   U1237 : NOR2_X1 port map( A1 => net92255, A2 => ALU_OPCODE(1), ZN => n252);
   U1154 : NOR2_X1 port map( A1 => net77056, A2 => net82508, ZN => n254);
   U256 : AOI21_X1 port map( B1 => n252, B2 => net77027, A => n254, ZN => n249)
                           ;
   U278 : NOR2_X1 port map( A1 => net83085, A2 => n304, ZN => n297);
   U280 : OAI21_X1 port map( B1 => net76624, B2 => net82650, A => n308, ZN => 
                           n307);
   U289 : NAND2_X1 port map( A1 => N2011, A2 => n320, ZN => n318);
   U1251 : NOR2_X1 port map( A1 => net77046, A2 => ALU_OPCODE(1), ZN => n1172);
   U1374 : NAND2_X1 port map( A1 => net92259, A2 => net74226, ZN => n1191);
   U1120 : NOR3_X1 port map( A1 => n1373, A2 => net92259, A3 => net76624, ZN =>
                           n1168);
   U1242 : NOR4_X1 port map( A1 => n1265, A2 => net74227, A3 => net92259, A4 =>
                           net82773, ZN => n1264);
   U277 : NOR3_X1 port map( A1 => net74226, A2 => net92259, A3 => net76624, ZN 
                           => n303);
   U276 : AOI21_X1 port map( B1 => net76624, B2 => n302, A => n303, ZN => n299)
                           ;
   U1287 : NOR2_X1 port map( A1 => net82508, A2 => net86253, ZN => n314);
   U1107 : AOI21_X1 port map( B1 => n301, B2 => net83925, A => net74253, ZN => 
                           n526);
   U1153 : AOI22_X1 port map( A1 => net92271, A2 => n1204, B1 => net83925, B2 
                           => n306, ZN => n1199);
   U275 : NAND2_X1 port map( A1 => net83925, A2 => n301, ZN => n300);
   U274 : OAI21_X1 port map( B1 => n299, B2 => net82639, A => n300, ZN => n298)
                           ;
   U273 : AOI22_X1 port map( A1 => n297, A2 => net92300, B1 => N2011, B2 => 
                           n298, ZN => n296);
   U272 : OAI21_X1 port map( B1 => n294, B2 => n295, A => n296, ZN => OVF);
   U357 : OAI21_X1 port map( B1 => n345, B2 => net82473, A => net76311, ZN => 
                           n427);
   U714 : OAI21_X1 port map( B1 => n345, B2 => DATA2(20), A => n1386, ZN => 
                           n828);
   U514 : AOI22_X1 port map( A1 => DATA1(28), A2 => n341, B1 => n1385, B2 => 
                           n1387, ZN => n630);
   U1051 : AOI21_X1 port map( B1 => net76297, B2 => net74295, A => net76555, ZN
                           => n1110);
   U916 : AOI21_X1 port map( B1 => n1385, B2 => net74386, A => net76555, ZN => 
                           n1005);
   U711 : OAI21_X1 port map( B1 => net76555, B2 => n830, A => DATA2(20), ZN => 
                           n829);
   U513 : NAND2_X1 port map( A1 => n630, A2 => net76311, ZN => n629);
   U512 : AOI22_X1 port map( A1 => n628, A2 => n519, B1 => DATA2(28), B2 => 
                           n629, ZN => n622);
   U1210 : NOR2_X1 port map( A1 => net83941, A2 => net74233, ZN => n1238);
   U1209 : NAND2_X1 port map( A1 => n1238, A2 => n315, ZN => n1237);
   U932 : AOI22_X1 port map( A1 => n1021, A2 => n508, B1 => DATA1(10), B2 => 
                           n1022, ZN => n1020);
   U1208 : OAI21_X1 port map( B1 => net82639, B2 => n1236, A => n1237, ZN => 
                           n508);
   U1243 : AOI21_X1 port map( B1 => net83941, B2 => net86253, A => net83927, ZN
                           => n1206);
   U1225 : NOR2_X1 port map( A1 => net83927, A2 => n314, ZN => n1253);
   U281 : AOI22_X1 port map( A1 => n309, A2 => n310, B1 => net92254, B2 => 
                           net83927, ZN => n308);
   U1361 : AOI22_X1 port map( A1 => n1274, A2 => n251, B1 => net83927, B2 => 
                           n1277, ZN => n1295);
   U1253 : AOI22_X1 port map( A1 => n310, A2 => n1273, B1 => n1274, B2 => 
                           net83927, ZN => n1272);
   U1118 : OAI21_X1 port map( B1 => net83941, B2 => net74228, A => net74224, ZN
                           => n1170);
   U1227 : NOR2_X1 port map( A1 => net77046, A2 => net74249, ZN => n1155);
   U1169 : OAI21_X1 port map( B1 => net74249, B2 => n1095, A => n1213, ZN => 
                           n582);
   U1033 : OAI33_X1 port map( A1 => n1094, A2 => net76732, A3 => net82639, B1 
                           => n1095, B2 => net76732, B3 => net74249, ZN => n352
                           );
   U1215 : NOR2_X1 port map( A1 => net74228, A2 => net74249, ZN => n1244);
   U1241 : AOI21_X1 port map( B1 => n1263, B2 => net82381, A => n1264, ZN => 
                           n1262);
   U1109 : OAI21_X1 port map( B1 => net74222, B2 => net74229, A => n1158, ZN =>
                           n1156);
   U1095 : OAI21_X1 port map( B1 => net82639, B2 => net74236, A => n1143, ZN =>
                           n350);
   U1368 : NOR4_X1 port map( A1 => net92259, A2 => net86253, A3 => net74222, A4
                           => net82639, ZN => n1338);
   U1367 : NOR2_X1 port map( A1 => n1208, A2 => n1338, ZN => n363);
   U1144 : OAI21_X1 port map( B1 => net76617, B2 => n289, A => n1193, ZN => 
                           CARRY);
   U929 : OAI21_X1 port map( B1 => net76617, B2 => n292, A => n1016, ZN => 
                           OUTALU(10));
   U660 : OAI21_X1 port map( B1 => net76617, B2 => n264, A => n782, ZN => 
                           OUTALU(20));
   U2 : OR2_X1 port map( A1 => n1171, A2 => net88905, ZN => n1173);
   U4 : NAND2_X1 port map( A1 => n1194, A2 => n1167, ZN => n1164);
   U6 : OR2_X1 port map( A1 => n1166, A2 => net88905, ZN => n1194);
   U11 : NOR2_X1 port map( A1 => DATA1(31), A2 => net82508, ZN => n1196);
   U12 : NOR2_X1 port map( A1 => N2010, A2 => n1341, ZN => n1198);
   U13 : OR2_X1 port map( A1 => n1198, A2 => n1340, ZN => n1354);
   U15 : OR2_X1 port map( A1 => net82508, A2 => n1348, ZN => n1341);
   U17 : INV_X1 port map( A => DATA1(31), ZN => net74284);
   U19 : NOR2_X1 port map( A1 => net83207, A2 => n1627_port, ZN => n1343);
   U20 : INV_X1 port map( A => n731, ZN => n1344);
   U21 : OR2_X1 port map( A1 => n1343, A2 => n1344, ZN => n1345);
   U23 : NOR2_X1 port map( A1 => n1343, A2 => n729, ZN => n1346);
   U25 : INV_X1 port map( A => net83955, ZN => n1348);
   U26 : NAND2_X1 port map( A1 => n1349, A2 => n1350, ZN => n294);
   U27 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n1349);
   U29 : NAND2_X1 port map( A1 => n1397, A2 => n1354, ZN => n1352);
   U30 : NAND2_X1 port map( A1 => n1352, A2 => n1353, ZN => n1350);
   U31 : OR2_X1 port map( A1 => n1348, A2 => net82650, ZN => n1353);
   U32 : NOR2_X1 port map( A1 => n1781, A2 => n1356, ZN => n1355);
   U33 : NAND2_X1 port map( A1 => n1384, A2 => n697, ZN => n1356);
   U37 : INV_X1 port map( A => n1359, ZN => n736);
   U42 : NOR2_X1 port map( A1 => n1345, A2 => n729, ZN => n1364);
   U44 : INV_X1 port map( A => N2008, ZN => n1367);
   U45 : NOR2_X1 port map( A1 => net83207, A2 => n1367, ZN => n1365);
   U47 : NAND2_X1 port map( A1 => n1369, A2 => n1370, ZN => n271);
   U48 : NAND2_X1 port map( A1 => N1639, A2 => net76327, ZN => n1369);
   U49 : NOR2_X1 port map( A1 => n1365, A2 => net82890, ZN => n1370);
   U52 : INV_X1 port map( A => n509, ZN => n1373);
   U54 : NOR2_X1 port map( A1 => n1373, A2 => net74248, ZN => n1371);
   U55 : INV_X1 port map( A => net82307, ZN => n1376);
   U56 : NAND2_X1 port map( A1 => n1377, A2 => n1378, ZN => n505);
   U57 : NAND2_X1 port map( A1 => N1641, A2 => net76329, ZN => n1377);
   U58 : NOR2_X1 port map( A1 => n1371, A2 => n1376, ZN => n1378);
   U59 : OAI21_X1 port map( B1 => net82819, B2 => n363, A => net82880, ZN => 
                           OUTALU(30));
   U65 : INV_X1 port map( A => n363, ZN => net74246);
   U66 : CLKBUF_X1 port map( A => net74246, Z => net76321);
   U68 : NOR2_X1 port map( A1 => n505, A2 => net82835, ZN => net82819);
   U72 : CLKBUF_X1 port map( A => n363, Z => net76617);
   U74 : INV_X1 port map( A => net92271, ZN => net82639);
   U75 : INV_X1 port map( A => n320, ZN => net74222);
   U77 : CLKBUF_X1 port map( A => ALU_OPCODE(4), Z => net86253);
   U78 : INV_X1 port map( A => net86253, ZN => net74226);
   U79 : NAND2_X1 port map( A1 => net92259, A2 => net86253, ZN => net82650);
   U87 : CLKBUF_X1 port map( A => n1772, Z => net76327);
   U89 : CLKBUF_X1 port map( A => n1772, Z => net76325);
   U90 : CLKBUF_X1 port map( A => n1772, Z => net76329);
   U91 : CLKBUF_X1 port map( A => n1172, Z => net82381);
   U92 : INV_X1 port map( A => n315, ZN => net74249);
   U93 : INV_X1 port map( A => net83927, ZN => net74228);
   U95 : CLKBUF_X1 port map( A => net86262, Z => net83927);
   U96 : NAND2_X1 port map( A1 => net88949, A2 => n1774, ZN => n503);
   U97 : OR2_X1 port map( A1 => net82639, A2 => n506, ZN => net82307);
   U98 : NAND2_X1 port map( A1 => n1420, A2 => net82307, ZN => net82867);
   U99 : AOI22_X1 port map( A1 => N1641, A2 => net76327, B1 => n508, B2 => n509
                           , ZN => net82949);
   U100 : INV_X1 port map( A => n508, ZN => net74248);
   U102 : NAND2_X1 port map( A1 => n1364, A2 => n717, ZN => n1381);
   U106 : OR2_X1 port map( A1 => n1425, A2 => n1427, ZN => n1383);
   U107 : OR2_X1 port map( A1 => net83207, A2 => n1626_port, ZN => n1384);
   U108 : NOR3_X1 port map( A1 => n271, A2 => n273, A3 => n1393, ZN => n270);
   U110 : NAND2_X1 port map( A1 => n1394, A2 => n620, ZN => n1393);
   U111 : NOR2_X1 port map( A1 => n1391, A2 => n274, ZN => n1394);
   U113 : INV_X1 port map( A => n1391, ZN => n1392);
   U114 : NAND2_X1 port map( A1 => n620, A2 => n1392, ZN => n272);
   U119 : INV_X1 port map( A => n488, ZN => n1386);
   U120 : CLKBUF_X1 port map( A => n1386, Z => net76311);
   U122 : INV_X1 port map( A => DATA1(28), ZN => n1387);
   U127 : INV_X1 port map( A => n345, ZN => n1385);
   U128 : CLKBUF_X1 port map( A => n1385, Z => net76297);
   U132 : AOI22_X1 port map( A1 => N1639, A2 => net76327, B1 => N2008, B2 => 
                           n362, ZN => net83203);
   U138 : NOR2_X1 port map( A1 => net82508, A2 => net82650, ZN => net83925);
   U140 : CLKBUF_X1 port map( A => ALU_OPCODE(5), Z => net82733);
   U141 : CLKBUF_X1 port map( A => ALU_OPCODE(6), Z => net76624);
   U143 : OR2_X1 port map( A1 => net92259, A2 => net86253, ZN => net83955);
   U145 : CLKBUF_X1 port map( A => ALU_OPCODE(1), Z => net92259);
   U146 : NOR2_X1 port map( A1 => net92255, A2 => net92259, ZN => net92254);
   U152 : NAND2_X1 port map( A1 => net92300, A2 => net83880, ZN => n317);
   U153 : OR2_X1 port map( A1 => n321, A2 => net82650, ZN => net83880);
   U157 : NOR2_X1 port map( A1 => ALU_OPCODE(5), A2 => net74226, ZN => net77027
                           );
   U160 : NOR2_X1 port map( A1 => n1414, A2 => net83085, ZN => net92271);
   U162 : INV_X1 port map( A => ALU_OPCODE(6), ZN => net92255);
   U169 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => net87788);
   U171 : NAND2_X1 port map( A1 => ALU_OPCODE(4), A2 => ALU_OPCODE(1), ZN => 
                           net77056);
   U174 : NAND2_X1 port map( A1 => N2010, A2 => n1165, ZN => n506);
   U175 : INV_X1 port map( A => N2010, ZN => net88905);
   U176 : NAND2_X1 port map( A1 => N2011, A2 => net87741, ZN => net87738);
   U177 : NAND2_X1 port map( A1 => N2011, A2 => net83893, ZN => net83237);
   U182 : OR2_X1 port map( A1 => net88905, A2 => net83853, ZN => net88949);
   U183 : NOR2_X1 port map( A1 => DATA1(31), A2 => DATA2(31), ZN => net88934);
   U184 : CLKBUF_X1 port map( A => DATA2(3), Z => n1403);
   U186 : INV_X1 port map( A => n1764, ZN => n1404);
   U190 : CLKBUF_X1 port map( A => DATA1(1), Z => n1405);
   U192 : OR2_X1 port map( A1 => net76617, A2 => n1795, ZN => n1407);
   U197 : NOR3_X1 port map( A1 => n1359, A2 => n275, A3 => n1595, ZN => n1409);
   U201 : OR2_X1 port map( A1 => n741, A2 => n1784, ZN => n1595);
   U206 : OR2_X1 port map( A1 => ALU_OPCODE(0), A2 => ALU_OPCODE(2), ZN => 
                           n1414);
   U210 : INV_X1 port map( A => net92254, ZN => net74235);
   U211 : OR2_X1 port map( A1 => n289, A2 => net76321, ZN => n1415);
   U212 : NAND2_X1 port map( A1 => net87738, A2 => n1401, ZN => n288);
   U213 : CLKBUF_X1 port map( A => DATA2(9), Z => n1416);
   U216 : NOR2_X1 port map( A1 => n1437, A2 => n1787, ZN => n1418);
   U217 : CLKBUF_X1 port map( A => net92255, Z => net83941);
   U218 : OR2_X1 port map( A1 => ALU_OPCODE(0), A2 => ALU_OPCODE(2), ZN => 
                           net83926);
   U220 : OR2_X1 port map( A1 => net83238, A2 => n1424, ZN => net83893);
   U221 : INV_X1 port map( A => n1199, ZN => net83238);
   U222 : INV_X1 port map( A => n1200, ZN => n1424);
   U225 : NOR2_X1 port map( A1 => n502, A2 => n504, ZN => n1420);
   U226 : OR2_X1 port map( A1 => n1421, A2 => n503, ZN => net82835);
   U227 : INV_X1 port map( A => n1420, ZN => n1421);
   U228 : NOR2_X1 port map( A1 => net83851, A2 => n1422, ZN => net83853);
   U229 : INV_X1 port map( A => n526, ZN => net83851);
   U230 : INV_X1 port map( A => n527, ZN => n1422);
   U232 : INV_X1 port map( A => n1208, ZN => net74233);
   U234 : INV_X1 port map( A => n1176, ZN => net74426);
   U236 : NOR2_X1 port map( A1 => n1426, A2 => net83207, ZN => n1427);
   U237 : INV_X1 port map( A => N2005, ZN => n1426);
   U238 : INV_X1 port map( A => n362, ZN => net83207);
   U240 : NAND2_X1 port map( A1 => net83203, A2 => net82891, ZN => n1429);
   U241 : AOI22_X1 port map( A1 => N1640, A2 => net76327, B1 => N2009, B2 => 
                           n362, ZN => n1430);
   U243 : CLKBUF_X1 port map( A => net74252, Z => net83091);
   U245 : CLKBUF_X1 port map( A => DATA2(12), Z => net83048);
   U248 : CLKBUF_X1 port map( A => DATA2(10), Z => n1432);
   U251 : NAND2_X1 port map( A1 => n646, A2 => n1780, ZN => n273);
   U253 : NOR2_X1 port map( A1 => n1436, A2 => net83207, ZN => n1437);
   U254 : INV_X1 port map( A => N2006, ZN => n1436);
   U261 : CLKBUF_X1 port map( A => DATA2(14), Z => n1438);
   U264 : NOR2_X1 port map( A1 => n1459, A2 => n1462, ZN => n1440);
   U268 : INV_X1 port map( A => net82890, ZN => net82891);
   U287 : NAND2_X1 port map( A1 => net83237, A2 => n1795, ZN => n1467);
   U423 : CLKBUF_X1 port map( A => ALU_OPCODE(2), Z => net82773);
   U435 : CLKBUF_X1 port map( A => DATA2(13), Z => n1448);
   U486 : CLKBUF_X1 port map( A => DATA2(11), Z => n1450);
   U504 : NOR2_X1 port map( A1 => n747, A2 => n1452, ZN => n1453);
   U525 : INV_X1 port map( A => n524, ZN => n1452);
   U604 : CLKBUF_X1 port map( A => DATA2(5), Z => n1456);
   U605 : CLKBUF_X1 port map( A => DATA2(6), Z => net82473);
   U638 : CLKBUF_X1 port map( A => DATA2(7), Z => n1457);
   U1163 : NAND2_X1 port map( A1 => n1466, A2 => n278, ZN => n1459);
   U1279 : CLKBUF_X1 port map( A => DATA2(8), Z => n1460);
   U1370 : NAND2_X1 port map( A1 => n1430, A2 => n1463, ZN => n284);
   U1375 : INV_X1 port map( A => n1462, ZN => n1463);
   U1376 : CLKBUF_X1 port map( A => DATA2(15), Z => n1464);
   U1381 : CLKBUF_X1 port map( A => n352, Z => net82287);
   U1382 : NOR3_X1 port map( A1 => n282, A2 => n283, A3 => n1606, ZN => n1466);
   U1383 : INV_X1 port map( A => net83926, ZN => n306);
   U1385 : INV_X1 port map( A => n1195, ZN => n1468);
   U1391 : INV_X1 port map( A => n411, ZN => n1618_port);
   U1392 : INV_X1 port map( A => n661, ZN => n1621_port);
   U1393 : INV_X1 port map( A => n534, ZN => n1674);
   U1394 : INV_X1 port map( A => n1551, ZN => n1673);
   U1396 : INV_X1 port map( A => n628, ZN => net74365);
   U1397 : INV_X1 port map( A => n359, ZN => n1662);
   U1402 : INV_X1 port map( A => n405, ZN => n1675);
   U1403 : INV_X1 port map( A => n456, ZN => n1664);
   U1404 : INV_X1 port map( A => n964, ZN => n1657);
   U1405 : INV_X1 port map( A => n415, ZN => n1656);
   U1406 : INV_X1 port map( A => n650, ZN => n1611_port);
   U1407 : INV_X1 port map( A => n333, ZN => n1652);
   U1408 : INV_X1 port map( A => n492, ZN => n1655);
   U1409 : INV_X1 port map( A => n361, ZN => n1672);
   U1410 : INV_X1 port map( A => n344, ZN => n1612_port);
   U1411 : INV_X1 port map( A => n658, ZN => n1663);
   U1412 : INV_X1 port map( A => n445, ZN => n1658);
   U1413 : CLKBUF_X1 port map( A => n514, Z => n1551);
   U1414 : INV_X1 port map( A => n519, ZN => net74293);
   U1418 : INV_X1 port map( A => n578, ZN => n1732);
   U1419 : INV_X1 port map( A => n462, ZN => n1736);
   U1420 : INV_X1 port map( A => n397, ZN => n1668);
   U1421 : CLKBUF_X1 port map( A => n1561, Z => n1475);
   U1423 : CLKBUF_X1 port map( A => n1568_port, Z => n1481);
   U1437 : INV_X1 port map( A => n563, ZN => n1679);
   U1438 : INV_X1 port map( A => n388, ZN => n1665);
   U1439 : INV_X1 port map( A => n601, ZN => n1610_port);
   U1440 : INV_X1 port map( A => n564, ZN => n1683);
   U1441 : INV_X1 port map( A => n819, ZN => n1681);
   U1442 : INV_X1 port map( A => n684, ZN => n1689);
   U1443 : INV_X1 port map( A => n356, ZN => n1669);
   U1444 : INV_X1 port map( A => n614, ZN => n1680);
   U1445 : INV_X1 port map( A => n407, ZN => n1687);
   U1446 : INV_X1 port map( A => n436, ZN => n1686);
   U1447 : INV_X1 port map( A => n419, ZN => n1678);
   U1448 : INV_X1 port map( A => n324, ZN => n1609);
   U1449 : INV_X1 port map( A => n941, ZN => n1598);
   U1450 : INV_X1 port map( A => n966, ZN => n1597);
   U1451 : INV_X1 port map( A => n894, ZN => n1600);
   U1452 : INV_X1 port map( A => n915, ZN => n1599);
   U1453 : INV_X1 port map( A => N1576, ZN => net74464);
   U1454 : INV_X1 port map( A => n1029, ZN => n1690);
   U1455 : INV_X1 port map( A => n510, ZN => n1768);
   U1460 : INV_X1 port map( A => n546, ZN => n1622_port);
   U1462 : INV_X1 port map( A => n1472, ZN => n1568_port);
   U1463 : INV_X1 port map( A => n428, ZN => n1701);
   U1464 : INV_X1 port map( A => n465, ZN => n1696);
   U1465 : INV_X1 port map( A => n1535, ZN => n1693);
   U1468 : INV_X1 port map( A => n747, ZN => n1671);
   U1469 : INV_X1 port map( A => n562, ZN => n1688);
   U1470 : INV_X1 port map( A => n522, ZN => n1670);
   U1471 : CLKBUF_X1 port map( A => n512, Z => n1555);
   U1472 : INV_X1 port map( A => n350, ZN => net74247);
   U1473 : INV_X1 port map( A => n703, ZN => n1667);
   U1476 : INV_X1 port map( A => n1126, ZN => n1661);
   U1477 : CLKBUF_X1 port map( A => n563, Z => n1538);
   U1478 : CLKBUF_X1 port map( A => n488, Z => net76555);
   U1479 : INV_X1 port map( A => n418, ZN => n1660);
   U1480 : CLKBUF_X1 port map( A => n341, Z => net76217);
   U1481 : INV_X1 port map( A => n713, ZN => n1666);
   U1484 : INV_X1 port map( A => n652, ZN => n1735);
   U1486 : INV_X1 port map( A => n781, ZN => n1731);
   U1487 : INV_X1 port map( A => n723, ZN => n1733);
   U1488 : CLKBUF_X1 port map( A => n356, Z => n1549);
   U1489 : CLKBUF_X1 port map( A => n357, Z => n1545);
   U1490 : INV_X1 port map( A => n408, ZN => n1717);
   U1493 : INV_X1 port map( A => n336, ZN => n1700);
   U1494 : INV_X1 port map( A => n285, ZN => n1606);
   U1495 : INV_X1 port map( A => n774, ZN => n1722);
   U1496 : INV_X1 port map( A => n1068, ZN => n1734);
   U1497 : INV_X1 port map( A => n473, ZN => n1713);
   U1499 : INV_X1 port map( A => n1145, ZN => net74236);
   U1502 : INV_X1 port map( A => n659, ZN => n1720);
   U1503 : INV_X1 port map( A => n639, ZN => n1710);
   U1505 : INV_X1 port map( A => n635, ZN => n1699);
   U1506 : INV_X1 port map( A => n682, ZN => n1724);
   U1507 : INV_X1 port map( A => n346, ZN => n1726);
   U1508 : INV_X1 port map( A => n1027, ZN => n1620_port);
   U1509 : INV_X1 port map( A => n1182, ZN => n1617_port);
   U1510 : INV_X1 port map( A => n808, ZN => n1682);
   U1511 : INV_X1 port map( A => n435, ZN => n1729);
   U1512 : INV_X1 port map( A => n1063, ZN => n1651);
   U1513 : INV_X1 port map( A => n530, ZN => n1730);
   U1514 : INV_X1 port map( A => n292, ZN => net74444);
   U1515 : INV_X1 port map( A => n281, ZN => n1608);
   U1516 : OR2_X1 port map( A1 => n1645, A2 => n510, ZN => n1470);
   U1517 : INV_X1 port map( A => n998, ZN => n1619_port);
   U1518 : INV_X1 port map( A => n983, ZN => n1613_port);
   U1519 : INV_X1 port map( A => n264, ZN => net74450);
   U1520 : INV_X1 port map( A => n1236, ZN => net74234);
   U1521 : INV_X1 port map( A => n827, ZN => n1635_port);
   U1522 : INV_X1 port map( A => N1999, ZN => n1634_port);
   U1523 : INV_X1 port map( A => N1577, ZN => net74463);
   U1524 : INV_X1 port map( A => n1251, ZN => n1588);
   U1525 : INV_X1 port map( A => N1572, ZN => n1589);
   U1526 : INV_X1 port map( A => net82287, ZN => net74362);
   U1527 : INV_X1 port map( A => net76732, ZN => net74367);
   U1528 : INV_X1 port map( A => n724, ZN => n1695);
   U1529 : INV_X1 port map( A => n370, ZN => n1614_port);
   U1530 : INV_X1 port map( A => n1181, ZN => n1641_port);
   U1531 : INV_X1 port map( A => n735, ZN => n1705);
   U1532 : INV_X1 port map( A => DATA1(16), ZN => n1752);
   U1533 : INV_X1 port map( A => DATA1(17), ZN => n1751);
   U1534 : INV_X1 port map( A => DATA1(9), ZN => n1758);
   U1535 : INV_X1 port map( A => DATA1(26), ZN => n1743);
   U1536 : INV_X1 port map( A => DATA1(27), ZN => n1742);
   U1537 : INV_X1 port map( A => DATA1(11), ZN => n1757);
   U1538 : INV_X1 port map( A => DATA1(10), ZN => net74264);
   U1539 : CLKBUF_X1 port map( A => n576, Z => n1535);
   U1540 : INV_X1 port map( A => n905, ZN => n1676);
   U1541 : INV_X1 port map( A => n582, ZN => net74250);
   U1542 : INV_X1 port map( A => n472, ZN => n1654);
   U1543 : CLKBUF_X1 port map( A => n465, Z => n1532);
   U1544 : INV_X1 port map( A => n387, ZN => n1691);
   U1546 : CLKBUF_X1 port map( A => n562, Z => n1540);
   U1547 : INV_X1 port map( A => n1405, ZN => n1766);
   U1549 : INV_X1 port map( A => n610, ZN => n1728);
   U1550 : INV_X1 port map( A => n251, ZN => net74229);
   U1551 : INV_X1 port map( A => n1179, ZN => n1624_port);
   U1555 : INV_X1 port map( A => n381, ZN => n1703);
   U1558 : INV_X1 port map( A => n926, ZN => n1718);
   U1559 : INV_X1 port map( A => n360, ZN => n1714);
   U1562 : INV_X1 port map( A => n800, ZN => n1727);
   U1564 : INV_X1 port map( A => n566, ZN => n1716);
   U1565 : INV_X1 port map( A => DATA1(6), ZN => n1761);
   U1566 : INV_X1 port map( A => DATA1(7), ZN => n1760);
   U1568 : INV_X1 port map( A => n438, ZN => n1723);
   U1569 : INV_X1 port map( A => n409, ZN => n1719);
   U1570 : INV_X1 port map( A => n460, ZN => n1715);
   U1571 : INV_X1 port map( A => n437, ZN => n1721);
   U1572 : INV_X1 port map( A => n498, ZN => n1706);
   U1573 : INV_X1 port map( A => n839, ZN => n1704);
   U1574 : INV_X1 port map( A => n376, ZN => n1708);
   U1575 : INV_X1 port map( A => DATA1(30), ZN => n1740);
   U1576 : INV_X1 port map( A => n1180, ZN => n1659);
   U1577 : INV_X1 port map( A => n491, ZN => n1707);
   U1578 : INV_X1 port map( A => n374, ZN => n1702);
   U1579 : INV_X1 port map( A => n725, ZN => n1711);
   U1580 : INV_X1 port map( A => n611, ZN => n1725);
   U1581 : INV_X1 port map( A => n301, ZN => net74243);
   U1582 : INV_X1 port map( A => n733, ZN => n1712);
   U1583 : INV_X1 port map( A => n547, ZN => n1684);
   U1584 : INV_X1 port map( A => n261, ZN => n1601);
   U1585 : INV_X1 port map( A => n751, ZN => n1694);
   U1586 : INV_X1 port map( A => n283, ZN => n1605);
   U1587 : INV_X1 port map( A => DATA1(14), ZN => n1754);
   U1588 : INV_X1 port map( A => DATA1(15), ZN => n1753);
   U1589 : INV_X1 port map( A => N1979, ZN => n1737);
   U1590 : INV_X1 port map( A => DATA1(5), ZN => n1762);
   U1591 : INV_X1 port map( A => DATA1(19), ZN => n1749);
   U1592 : INV_X1 port map( A => n1289, ZN => n1629_port);
   U1593 : INV_X1 port map( A => n636, ZN => n1709);
   U1594 : INV_X1 port map( A => n486, ZN => n1677);
   U1595 : INV_X1 port map( A => n332, ZN => n1653);
   U1596 : INV_X1 port map( A => n1112, ZN => n1770);
   U1597 : INV_X1 port map( A => N2003, ZN => n1627_port);
   U1598 : INV_X1 port map( A => N1998, ZN => n1636_port);
   U1599 : INV_X1 port map( A => N1995, ZN => n1644);
   U1600 : INV_X1 port map( A => N1997, ZN => n1639_port);
   U1601 : INV_X1 port map( A => N1996, ZN => n1642);
   U1602 : INV_X1 port map( A => N2000, ZN => n1633_port);
   U1603 : INV_X1 port map( A => N2004, ZN => n1626_port);
   U1604 : INV_X1 port map( A => N2002, ZN => n1631_port);
   U1605 : INV_X1 port map( A => N2001, ZN => n1632_port);
   U1620 : INV_X1 port map( A => n1306, ZN => n1637_port);
   U1621 : INV_X1 port map( A => n1154, ZN => net74253);
   U1622 : INV_X1 port map( A => n1336, ZN => n1625_port);
   U1623 : INV_X1 port map( A => n1178, ZN => n1630_port);
   U1624 : INV_X1 port map( A => DATA1(21), ZN => n1748);
   U1625 : INV_X1 port map( A => DATA1(25), ZN => n1744);
   U1626 : INV_X1 port map( A => DATA1(8), ZN => n1759);
   U1627 : INV_X1 port map( A => n496, ZN => n1685);
   U1628 : INV_X1 port map( A => n425, ZN => n1615_port);
   U1629 : INV_X1 port map( A => n393, ZN => n1616_port);
   U1632 : INV_X1 port map( A => n485, ZN => n1697);
   U1639 : INV_X1 port map( A => n1275, ZN => n1739);
   U1640 : CLKBUF_X1 port map( A => DATA2(4), Z => net76732);
   U1641 : INV_X1 port map( A => n1403, ZN => n1692);
   U1643 : INV_X1 port map( A => DATA2(1), ZN => net74295);
   U1644 : INV_X1 port map( A => n310, ZN => net74225);
   U1645 : INV_X1 port map( A => DATA2(2), ZN => n1698);
   U1654 : INV_X1 port map( A => DATA1(4), ZN => n1763);
   U1655 : INV_X1 port map( A => n1461, ZN => n1765);
   U1657 : INV_X1 port map( A => DATA2(19), ZN => n1638_port);
   U1658 : INV_X1 port map( A => DATA1(12), ZN => n1756);
   U1660 : INV_X1 port map( A => DATA2(0), ZN => n1738);
   U1661 : INV_X1 port map( A => DATA1(13), ZN => n1755);
   U1662 : INV_X1 port map( A => DATA1(29), ZN => n1741);
   U1663 : INV_X1 port map( A => DATA1(24), ZN => n1745);
   U1664 : INV_X1 port map( A => DATA1(18), ZN => n1750);
   U1666 : INV_X1 port map( A => DATA1(22), ZN => n1747);
   U1667 : INV_X1 port map( A => DATA1(23), ZN => n1746);
   U1668 : INV_X1 port map( A => n1432, ZN => n1649);
   U1669 : OR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n1471);
   U1670 : OR2_X1 port map( A1 => net74295, A2 => DATA2(0), ZN => n1472);
   U1671 : INV_X1 port map( A => n829, ZN => net74400);
   U1672 : INV_X1 port map( A => n314, ZN => net74224);
   U1673 : INV_X1 port map( A => n1206, ZN => net74227);
   U1674 : INV_X1 port map( A => net83048, ZN => net74386);
   U1675 : INV_X1 port map( A => n1438, ZN => n1647);
   U1676 : INV_X1 port map( A => n1450, ZN => n1648);
   U1677 : INV_X1 port map( A => DATA2(16), ZN => n1645);
   U1678 : INV_X1 port map( A => DATA2(18), ZN => n1640_port);
   U1679 : INV_X1 port map( A => DATA2(24), ZN => n1628_port);
   U1680 : INV_X1 port map( A => n1416, ZN => n1650);
   U1681 : INV_X1 port map( A => DATA2(17), ZN => n1643);
   U1682 : INV_X1 port map( A => n506, ZN => net74455);
   U1683 : INV_X1 port map( A => n1429, ZN => n1604);
   U1684 : INV_X1 port map( A => n272, ZN => net74436);
   U1685 : INV_X1 port map( A => n619, ZN => OUTALU(27));
   U1686 : INV_X1 port map( A => n643, ZN => OUTALU(26));
   U1687 : INV_X1 port map( A => n876, ZN => OUTALU(16));
   U1688 : INV_X1 port map( A => n858, ZN => OUTALU(17));
   U1689 : INV_X1 port map( A => n822, ZN => OUTALU(19));
   U1690 : INV_X1 port map( A => n840, ZN => OUTALU(18));
   U1691 : INV_X1 port map( A => n801, ZN => OUTALU(1));
   U1692 : INV_X1 port map( A => n280, ZN => n1607);
   U1693 : INV_X1 port map( A => n1192, ZN => n1769);
   U1694 : INV_X1 port map( A => n1399, ZN => n1767);
   U1695 : INV_X1 port map( A => net92259, ZN => net74238);
   U1696 : AND2_X2 port map( A1 => ALU_OPCODE(2), A2 => net74252, ZN => n315);
   U1697 : INV_X1 port map( A => ALU_OPCODE(0), ZN => net74252);
   U1698 : INV_X1 port map( A => net82773, ZN => net74231);
   U1699 : INV_X1 port map( A => ALU_OPCODE(3), ZN => net77046);
   U1700 : INV_X1 port map( A => n1464, ZN => n1646);
   U1712 : INV_X1 port map( A => n520, ZN => n1577_port);
   U1715 : INV_X1 port map( A => n518, ZN => n1585);
   r167 : ALU_N32_DW01_cmp6_0 port map( A(31) => DATA1(31), A(30) => DATA1(30),
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => n1404, A(2) => n1461, A(1) => 
                           n1405, A(0) => n1399, B(31) => DATA2(31), B(30) => 
                           DATA2(30), B(29) => DATA2(29), B(28) => DATA2(28), 
                           B(27) => DATA2(27), B(26) => DATA2(26), B(25) => 
                           DATA2(25), B(24) => DATA2(24), B(23) => DATA2(23), 
                           B(22) => DATA2(22), B(21) => DATA2(21), B(20) => 
                           DATA2(20), B(19) => DATA2(19), B(18) => DATA2(18), 
                           B(17) => DATA2(17), B(16) => DATA2(16), B(15) => 
                           n1464, B(14) => n1438, B(13) => n1448, B(12) => 
                           net83048, B(11) => n1450, B(10) => n1432, B(9) => 
                           n1416, B(8) => n1460, B(7) => n1457, B(6) => 
                           net82473, B(5) => n1456, B(4) => net76732, B(3) => 
                           n1403, B(2) => DATA2(2), B(1) => DATA2(1), B(0) => 
                           DATA2(0), TC => n3, LT => n_1065, GT => n_1066, EQ 
                           => n_1067, LE => N1572, GE => N1573, NE => n_1068);
   r166 : ALU_N32_DW01_cmp6_1 port map( A(31) => DATA1(31), A(30) => DATA1(30),
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => n1404, A(2) => n1461, A(1) => 
                           n1405, A(0) => n1399, B(31) => DATA2(31), B(30) => 
                           DATA2(30), B(29) => DATA2(29), B(28) => DATA2(28), 
                           B(27) => DATA2(27), B(26) => DATA2(26), B(25) => 
                           DATA2(25), B(24) => DATA2(24), B(23) => DATA2(23), 
                           B(22) => DATA2(22), B(21) => DATA2(21), B(20) => 
                           DATA2(20), B(19) => DATA2(19), B(18) => DATA2(18), 
                           B(17) => DATA2(17), B(16) => DATA2(16), B(15) => 
                           n1464, B(14) => n1438, B(13) => n1448, B(12) => 
                           net83048, B(11) => n1450, B(10) => n1432, B(9) => 
                           n1416, B(8) => n1460, B(7) => n1457, B(6) => 
                           net82473, B(5) => n1456, B(4) => net76732, B(3) => 
                           n1403, B(2) => DATA2(2), B(1) => DATA2(1), B(0) => 
                           DATA2(0), TC => n4, LT => n_1069, GT => n_1070, EQ 
                           => N1568, LE => N1576, GE => N1577, NE => n_1071);
   r79 : ALU_N32_DW02_mult_0 port map( A(15) => DATA1(15), A(14) => DATA1(14), 
                           A(13) => DATA1(13), A(12) => DATA1(12), A(11) => 
                           DATA1(11), A(10) => DATA1(10), A(9) => DATA1(9), 
                           A(8) => DATA1(8), A(7) => DATA1(7), A(6) => DATA1(6)
                           , A(5) => DATA1(5), A(4) => DATA1(4), A(3) => 
                           DATA1(3), A(2) => DATA1(2), A(1) => DATA1(1), A(0) 
                           => DATA1(0), B(15) => DATA2(15), B(14) => DATA2(14),
                           B(13) => DATA2(13), B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6)
                           , B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), TC => U2_U1_Z_0, PRODUCT(31) => N1641, 
                           PRODUCT(30) => N1640, PRODUCT(29) => N1639, 
                           PRODUCT(28) => N1638, PRODUCT(27) => N1637, 
                           PRODUCT(26) => N1636, PRODUCT(25) => N1635, 
                           PRODUCT(24) => N1634, PRODUCT(23) => N1633, 
                           PRODUCT(22) => N1632, PRODUCT(21) => N1631, 
                           PRODUCT(20) => N1630, PRODUCT(19) => N1629, 
                           PRODUCT(18) => N1628, PRODUCT(17) => N1627, 
                           PRODUCT(16) => N1626, PRODUCT(15) => N1625, 
                           PRODUCT(14) => N1624, PRODUCT(13) => N1623, 
                           PRODUCT(12) => N1622, PRODUCT(11) => N1621, 
                           PRODUCT(10) => N1620, PRODUCT(9) => N1619, 
                           PRODUCT(8) => N1618, PRODUCT(7) => N1617, PRODUCT(6)
                           => N1616, PRODUCT(5) => N1615, PRODUCT(4) => N1614, 
                           PRODUCT(3) => N1613, PRODUCT(2) => N1612, PRODUCT(1)
                           => N1611, PRODUCT(0) => N1610);
   r170 : ALU_N32_DW01_addsub_3 port map( A(32) => n1, A(31) => DATA1(31), 
                           A(30) => DATA1(30), A(29) => DATA1(29), A(28) => 
                           DATA1(28), A(27) => DATA1(27), A(26) => DATA1(26), 
                           A(25) => DATA1(25), A(24) => DATA1(24), A(23) => 
                           DATA1(23), A(22) => DATA1(22), A(21) => DATA1(21), 
                           A(20) => DATA1(20), A(19) => DATA1(19), A(18) => 
                           DATA1(18), A(17) => DATA1(17), A(16) => DATA1(16), 
                           A(15) => DATA1(15), A(14) => DATA1(14), A(13) => 
                           DATA1(13), A(12) => DATA1(12), A(11) => DATA1(11), 
                           A(10) => DATA1(10), A(9) => DATA1(9), A(8) => 
                           DATA1(8), A(7) => DATA1(7), A(6) => DATA1(6), A(5) 
                           => DATA1(5), A(4) => DATA1(4), A(3) => n1404, A(2) 
                           => n1461, A(1) => n1405, A(0) => n1399, B(32) => n1,
                           B(31) => DATA2(31), B(30) => DATA2(30), B(29) => 
                           DATA2(29), B(28) => DATA2(28), B(27) => DATA2(27), 
                           B(26) => DATA2(26), B(25) => DATA2(25), B(24) => 
                           DATA2(24), B(23) => DATA2(23), B(22) => DATA2(22), 
                           B(21) => DATA2(21), B(20) => DATA2(20), B(19) => 
                           DATA2(19), B(18) => DATA2(18), B(17) => DATA2(17), 
                           B(16) => DATA2(16), B(15) => n1464, B(14) => n1438, 
                           B(13) => n1448, B(12) => net83048, B(11) => n1450, 
                           B(10) => n1432, B(9) => n1416, B(8) => n1460, B(7) 
                           => n1457, B(6) => net82473, B(5) => n1456, B(4) => 
                           DATA2(4), B(3) => n1403, B(2) => DATA2(2), B(1) => 
                           DATA2(1), B(0) => DATA2(0), CI => n2, ADD_SUB => 
                           n1339, SUM(32) => N2011, SUM(31) => N2010, SUM(30) 
                           => N2009, SUM(29) => N2008, SUM(28) => N2007, 
                           SUM(27) => N2006, SUM(26) => N2005, SUM(25) => N2004
                           , SUM(24) => N2003, SUM(23) => N2002, SUM(22) => 
                           N2001, SUM(21) => N2000, SUM(20) => N1999, SUM(19) 
                           => N1998, SUM(18) => N1997, SUM(17) => N1996, 
                           SUM(16) => N1995, SUM(15) => N1994, SUM(14) => N1993
                           , SUM(13) => N1992, SUM(12) => N1991, SUM(11) => 
                           N1990, SUM(10) => N1989, SUM(9) => N1988, SUM(8) => 
                           N1987, SUM(7) => N1986, SUM(6) => N1985, SUM(5) => 
                           N1984, SUM(4) => N1983, SUM(3) => N1982, SUM(2) => 
                           N1981, SUM(1) => N1980, SUM(0) => N1979, CO => 
                           n_1072);
   U3 : INV_X2 port map( A => ALU_OPCODE(5), ZN => net82508);
   U10 : AND2_X1 port map( A1 => net77050, A2 => n1474, ZN => U2_U1_Z_0);
   U14 : AND2_X1 port map( A1 => n321, A2 => net82381, ZN => n1771);
   U16 : AND2_X1 port map( A1 => N1641, A2 => n1771, ZN => n1357);
   U18 : AND2_X1 port map( A1 => n1244, A2 => net82381, ZN => n1772);
   U22 : AND2_X1 port map( A1 => n766, A2 => n767, ZN => n1773);
   U24 : NOR2_X1 port map( A1 => n1785, A2 => n1453, ZN => n1774);
   U28 : AND2_X1 port map( A1 => net87738, A2 => n1407, ZN => n1775);
   U34 : AND2_X1 port map( A1 => n259, A2 => n260, ZN => n1776);
   U35 : OR2_X1 port map( A1 => n1599, A2 => n1600, ZN => n1777);
   U36 : OR2_X1 port map( A1 => n1777, A2 => n288, ZN => n1778);
   U38 : OR4_X1 port map( A1 => DATA2(19), A2 => n1624_port, A3 => n1185, A4 =>
                           n1186, ZN => n1779);
   U39 : AND3_X1 port map( A1 => n647, A2 => n644, A3 => n645, ZN => n1780);
   U40 : OR3_X1 port map( A1 => n694, A2 => n693, A3 => n695, ZN => n1781);
   U41 : AND2_X1 port map( A1 => n778, A2 => n779, ZN => n1782);
   U43 : OR3_X1 port map( A1 => net74293, A2 => n1207, A3 => n1675, ZN => n1783
                           );
   U46 : OR3_X1 port map( A1 => n740, A2 => n738, A3 => n739, ZN => n1784);
   U50 : NOR2_X1 port map( A1 => n1730, A2 => n522, ZN => n1785);
   U51 : AND2_X1 port map( A1 => DATA2(31), A2 => DATA1(31), ZN => n1786);
   U53 : NOR2_X1 port map( A1 => n510, A2 => n1648, ZN => n1787);
   U60 : NAND2_X1 port map( A1 => n687, A2 => n1788, ZN => n274);
   U61 : NOR2_X1 port map( A1 => n1789, A2 => n1383, ZN => n1788);
   U62 : NOR2_X1 port map( A1 => n510, A2 => n1649, ZN => n1789);
   U63 : AND2_X1 port map( A1 => net82949, A2 => n1790, ZN => n287);
   U64 : NOR2_X1 port map( A1 => n1791, A2 => n1778, ZN => n1790);
   U67 : OR2_X1 port map( A1 => n503, A2 => net82867, ZN => n1791);
   U69 : NOR4_X2 port map( A1 => n783, A2 => n784, A3 => n785, A4 => n786, ZN 
                           => n264);
   U70 : AND2_X1 port map( A1 => n1377, A2 => n1792, ZN => net77055);
   U71 : AND2_X1 port map( A1 => n1378, A2 => n1793, ZN => n1792);
   U73 : INV_X1 port map( A => net82835, ZN => n1793);
   U76 : AND2_X1 port map( A1 => n1776, A2 => n286, ZN => n1794);
   U80 : AND3_X1 port map( A1 => net82699, A2 => n1447, A3 => n1794, ZN => 
                           n1465);
   U81 : NAND2_X1 port map( A1 => n284, A2 => net76617, ZN => net82880);
   U82 : INV_X1 port map( A => DATA1(3), ZN => n1764);
   U83 : AND2_X1 port map( A1 => n1346, A2 => n731, ZN => n716);
   U84 : AND2_X1 port map( A1 => net83893, A2 => net76321, ZN => net87741);
   U85 : AND2_X1 port map( A1 => net92255, A2 => n1172, ZN => n1474);
   U86 : AND2_X1 port map( A1 => net86262, A2 => n315, ZN => net77050);
   U88 : AND2_X1 port map( A1 => net83955, A2 => n1196, ZN => n1340);
   U94 : MUX2_X1 port map( A => N2010, B => DATA1(31), S => DATA2(31), Z => 
                           n1397);
   U101 : CLKBUF_X1 port map( A => DATA1(2), Z => n1461);
   U103 : CLKBUF_X1 port map( A => ALU_OPCODE(3), Z => net83085);
   U104 : AND2_X1 port map( A1 => n1415, A2 => n1407, ZN => n1401);
   U105 : AND2_X1 port map( A1 => n270, A2 => n269, ZN => net82699);
   U109 : AND2_X1 port map( A1 => n1409, A2 => n1355, ZN => n269);
   U112 : AND2_X1 port map( A1 => n1430, A2 => n1440, ZN => n1447);
   U115 : AND2_X1 port map( A1 => net82733, A2 => net86253, ZN => n251);
   U116 : AND2_X1 port map( A1 => net82508, A2 => ALU_OPCODE(4), ZN => net86262
                           );
   U117 : AND2_X1 port map( A1 => n592, A2 => n1549, ZN => n585);
   U118 : NAND4_X1 port map( A1 => n1285, A2 => n1286, A3 => n1287, A4 => n1288
                           , ZN => n1073);
   U121 : AND2_X1 port map( A1 => n1535, A2 => n776, ZN => n775);
   U123 : CLKBUF_X1 port map( A => DATA1(0), Z => n1399);
   U124 : AND2_X1 port map( A1 => n588, A2 => n361, ZN => n587);
   U125 : AND2_X1 port map( A1 => net87788, A2 => net92271, ZN => n1339);
   U126 : NAND3_X1 port map( A1 => n572, A2 => n570, A3 => n571, ZN => n1462);
   U129 : AND3_X1 port map( A1 => n1468, A2 => n1783, A3 => n1470, ZN => n1795)
                           ;
   U130 : INV_X1 port map( A => n1174, ZN => n1171);
   U131 : NOR2_X1 port map( A1 => n1796, A2 => n1797, ZN => n1157);
   U133 : OR3_X1 port map( A1 => net83091, A2 => net86253, A3 => n321, ZN => 
                           n1796);
   U134 : OR3_X1 port map( A1 => net83085, A2 => net82773, A3 => net92259, ZN 
                           => n1797);
   U135 : MUX2_X1 port map( A => n1786, B => net88934, S => N2010, Z => 
                           net92300);
   U136 : INV_X1 port map( A => n764, ZN => n1363);
   U137 : NAND3_X1 port map( A1 => n621, A2 => n623, A3 => n622, ZN => n1391);
   U139 : NAND3_X1 port map( A1 => n597, A2 => n599, A3 => n598, ZN => net82890
                           );
   U142 : NAND4_X1 port map( A1 => n802, A2 => n803, A3 => n804, A4 => n805, ZN
                           => n261);
   U144 : NAND4_X1 port map( A1 => n539, A2 => n540, A3 => n541, A4 => n542, ZN
                           => n283);
   U147 : NAND4_X1 port map( A1 => n478, A2 => n479, A3 => n480, A4 => n481, ZN
                           => n282);
   U148 : NAND4_X1 port map( A1 => n422, A2 => n423, A3 => n424, A4 => 
                           n1615_port, ZN => n280);
   U149 : NAND4_X1 port map( A1 => n390, A2 => n391, A3 => n392, A4 => 
                           n1616_port, ZN => n279);
   U150 : NAND4_X1 port map( A1 => n1017, A2 => n1018, A3 => n1019, A4 => n1020
                           , ZN => n291);
   U151 : NAND4_X1 port map( A1 => n1782, A2 => n1361, A3 => n1773, A4 => n1363
                           , ZN => n1359);
   U154 : INV_X1 port map( A => n762, ZN => n1361);
   U155 : NAND3_X1 port map( A1 => n673, A2 => n670, A3 => n671, ZN => n1425);
   U156 : AND2_X1 port map( A1 => n665, A2 => n1418, ZN => n646);
   U158 : AND2_X1 port map( A1 => n1465, A2 => n287, ZN => ZERO);
   U159 : INV_X2 port map( A => n1577_port, ZN => n1573_port);
   U161 : INV_X2 port map( A => n1585, ZN => n1582);
   U163 : INV_X2 port map( A => n1471, ZN => n1561);
   U164 : OAI21_X2 port map( B1 => n1153, B2 => net82639, A => n526, ZN => n362
                           );

end SYN_ARITH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_mux21_N32_3 is

   port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m : 
         out std_logic_vector (31 downto 0));

end gen_mux21_N32_3;

architecture SYN_dflow of gen_mux21_N32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63
      , n64, n65, n62, n66, n68, n70, n71, n73, n74, n75, n77, n81, n82, n83, 
      n84, n85, n86 : std_logic;

begin
   
   U34 : AOI22_X1 port map( A1 => x(9), A2 => n82, B1 => y(9), B2 => n86, ZN =>
                           n34);
   U35 : AOI22_X1 port map( A1 => x(8), A2 => n68, B1 => y(8), B2 => n86, ZN =>
                           n35);
   U36 : AOI22_X1 port map( A1 => x(7), A2 => n82, B1 => y(7), B2 => n86, ZN =>
                           n36);
   U37 : AOI22_X1 port map( A1 => x(6), A2 => n82, B1 => y(6), B2 => n77, ZN =>
                           n37);
   U38 : AOI22_X1 port map( A1 => x(5), A2 => n82, B1 => y(5), B2 => n77, ZN =>
                           n38);
   U39 : AOI22_X1 port map( A1 => x(4), A2 => n82, B1 => y(4), B2 => n77, ZN =>
                           n39);
   U40 : AOI22_X1 port map( A1 => x(3), A2 => n68, B1 => y(3), B2 => n86, ZN =>
                           n40);
   U41 : AOI22_X1 port map( A1 => x(31), A2 => n83, B1 => y(31), B2 => n75, ZN 
                           => n41);
   U42 : AOI22_X1 port map( A1 => x(30), A2 => n83, B1 => y(30), B2 => n75, ZN 
                           => n42);
   U43 : AOI22_X1 port map( A1 => x(2), A2 => n82, B1 => y(2), B2 => n86, ZN =>
                           n43);
   U44 : AOI22_X1 port map( A1 => x(29), A2 => n83, B1 => y(29), B2 => n75, ZN 
                           => n44);
   U45 : AOI22_X1 port map( A1 => x(28), A2 => n83, B1 => y(28), B2 => n75, ZN 
                           => n45);
   U46 : AOI22_X1 port map( A1 => x(27), A2 => n83, B1 => y(27), B2 => n75, ZN 
                           => n46);
   U47 : AOI22_X1 port map( A1 => x(26), A2 => n83, B1 => y(26), B2 => n75, ZN 
                           => n47);
   U48 : AOI22_X1 port map( A1 => x(25), A2 => n83, B1 => y(25), B2 => n75, ZN 
                           => n48);
   U49 : AOI22_X1 port map( A1 => x(24), A2 => n83, B1 => y(24), B2 => n75, ZN 
                           => n49);
   U50 : AOI22_X1 port map( A1 => x(23), A2 => n83, B1 => y(23), B2 => n75, ZN 
                           => n50);
   U51 : AOI22_X1 port map( A1 => x(22), A2 => n83, B1 => y(22), B2 => n75, ZN 
                           => n51);
   U52 : AOI22_X1 port map( A1 => x(21), A2 => n83, B1 => y(21), B2 => n75, ZN 
                           => n52);
   U53 : AOI22_X1 port map( A1 => x(20), A2 => n83, B1 => y(20), B2 => n75, ZN 
                           => n53);
   U54 : AOI22_X1 port map( A1 => n82, A2 => x(1), B1 => n86, B2 => y(1), ZN =>
                           n54);
   U55 : AOI22_X1 port map( A1 => x(19), A2 => n83, B1 => y(19), B2 => n75, ZN 
                           => n55);
   U56 : AOI22_X1 port map( A1 => x(18), A2 => n83, B1 => y(18), B2 => n75, ZN 
                           => n56);
   U57 : AOI22_X1 port map( A1 => x(17), A2 => n83, B1 => y(17), B2 => n75, ZN 
                           => n57);
   U58 : AOI22_X1 port map( A1 => x(16), A2 => n83, B1 => y(16), B2 => n75, ZN 
                           => n58);
   U59 : AOI22_X1 port map( A1 => n70, A2 => x(15), B1 => n73, B2 => y(15), ZN 
                           => n59);
   U60 : AOI22_X1 port map( A1 => n74, A2 => x(14), B1 => n71, B2 => y(14), ZN 
                           => n60);
   U61 : AOI22_X1 port map( A1 => n74, A2 => x(13), B1 => n71, B2 => y(13), ZN 
                           => n61);
   U63 : AOI22_X1 port map( A1 => n68, A2 => x(11), B1 => y(11), B2 => n85, ZN 
                           => n63);
   U64 : AOI22_X1 port map( A1 => x(10), A2 => n70, B1 => y(10), B2 => n81, ZN 
                           => n64);
   U65 : AOI22_X1 port map( A1 => n82, A2 => x(0), B1 => n73, B2 => y(0), ZN =>
                           n65);
   U2 : NAND2_X1 port map( A1 => n68, A2 => x(12), ZN => n62);
   U3 : NAND2_X1 port map( A1 => y(12), A2 => n85, ZN => n66);
   U4 : NAND2_X1 port map( A1 => n62, A2 => n66, ZN => m(12));
   U5 : INV_X1 port map( A => n81, ZN => n68);
   U12 : INV_X1 port map( A => n81, ZN => n70);
   U16 : INV_X1 port map( A => n75, ZN => n83);
   U17 : CLKBUF_X1 port map( A => n86, Z => n75);
   U18 : INV_X1 port map( A => n84, ZN => n74);
   U22 : INV_X1 port map( A => n64, ZN => m(10));
   U24 : INV_X1 port map( A => n54, ZN => m(1));
   U25 : INV_X1 port map( A => n60, ZN => m(14));
   U26 : INV_X1 port map( A => n34, ZN => m(9));
   U27 : INV_X1 port map( A => n61, ZN => m(13));
   U28 : INV_X1 port map( A => n63, ZN => m(11));
   U29 : INV_X1 port map( A => n40, ZN => m(3));
   U30 : INV_X1 port map( A => n38, ZN => m(5));
   U31 : INV_X1 port map( A => n43, ZN => m(2));
   U32 : INV_X1 port map( A => n35, ZN => m(8));
   U33 : INV_X1 port map( A => n36, ZN => m(7));
   U62 : INV_X1 port map( A => n37, ZN => m(6));
   U66 : INV_X1 port map( A => n39, ZN => m(4));
   U67 : INV_X1 port map( A => n65, ZN => m(0));
   U68 : INV_X1 port map( A => n52, ZN => m(21));
   U69 : INV_X1 port map( A => n53, ZN => m(20));
   U70 : INV_X1 port map( A => n55, ZN => m(19));
   U71 : INV_X1 port map( A => n57, ZN => m(17));
   U72 : INV_X1 port map( A => n58, ZN => m(16));
   U73 : INV_X1 port map( A => n56, ZN => m(18));
   U74 : INV_X1 port map( A => n51, ZN => m(22));
   U75 : INV_X1 port map( A => n44, ZN => m(29));
   U76 : INV_X1 port map( A => n42, ZN => m(30));
   U77 : INV_X1 port map( A => n46, ZN => m(27));
   U78 : INV_X1 port map( A => n45, ZN => m(28));
   U79 : INV_X1 port map( A => n48, ZN => m(25));
   U80 : INV_X1 port map( A => n47, ZN => m(26));
   U81 : INV_X1 port map( A => n41, ZN => m(31));
   U82 : INV_X1 port map( A => n50, ZN => m(23));
   U83 : INV_X1 port map( A => n49, ZN => m(24));
   U84 : INV_X1 port map( A => n59, ZN => m(15));
   U85 : INV_X1 port map( A => n71, ZN => n82);
   U1 : BUF_X1 port map( A => n73, Z => n77);
   U6 : BUF_X1 port map( A => n84, Z => n86);
   U7 : BUF_X1 port map( A => sel, Z => n84);
   U8 : BUF_X1 port map( A => sel, Z => n71);
   U9 : BUF_X1 port map( A => sel, Z => n81);
   U10 : BUF_X1 port map( A => n84, Z => n85);
   U11 : BUF_X1 port map( A => n71, Z => n73);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_mux21_N32_0 is

   port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m : 
         out std_logic_vector (31 downto 0));

end gen_mux21_N32_0;

architecture SYN_dflow of gen_mux21_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, net75115, net75113, net75109, net76536, net81028, net82506, 
      n33, n65, n67, n68 : std_logic;

begin
   
   U34 : AOI22_X1 port map( A1 => x(9), A2 => net76536, B1 => y(9), B2 => 
                           net75115, ZN => n34);
   U35 : AOI22_X1 port map( A1 => x(8), A2 => net75109, B1 => y(8), B2 => 
                           net75115, ZN => n35);
   U36 : AOI22_X1 port map( A1 => x(7), A2 => net76536, B1 => y(7), B2 => 
                           net75113, ZN => n36);
   U37 : AOI22_X1 port map( A1 => x(6), A2 => net75109, B1 => y(6), B2 => 
                           net75115, ZN => n37);
   U38 : AOI22_X1 port map( A1 => x(5), A2 => net76536, B1 => y(5), B2 => 
                           net75113, ZN => n38);
   U39 : AOI22_X1 port map( A1 => x(4), A2 => net76536, B1 => y(4), B2 => 
                           net75115, ZN => n39);
   U40 : AOI22_X1 port map( A1 => x(3), A2 => net76536, B1 => y(3), B2 => 
                           net75113, ZN => n40);
   U41 : AOI22_X1 port map( A1 => x(31), A2 => net75109, B1 => y(31), B2 => 
                           net75113, ZN => n41);
   U42 : AOI22_X1 port map( A1 => x(30), A2 => net76536, B1 => y(30), B2 => 
                           net75113, ZN => n42);
   U43 : AOI22_X1 port map( A1 => net81028, A2 => x(2), B1 => y(2), B2 => 
                           net82506, ZN => n43);
   U44 : AOI22_X1 port map( A1 => x(29), A2 => net76536, B1 => y(29), B2 => 
                           net75115, ZN => n44);
   U45 : AOI22_X1 port map( A1 => x(28), A2 => net75109, B1 => y(28), B2 => 
                           net75113, ZN => n45);
   U46 : AOI22_X1 port map( A1 => x(27), A2 => net75109, B1 => y(27), B2 => 
                           net75115, ZN => n46);
   U47 : AOI22_X1 port map( A1 => x(26), A2 => net75109, B1 => y(26), B2 => 
                           net75115, ZN => n47);
   U48 : AOI22_X1 port map( A1 => x(25), A2 => net75109, B1 => y(25), B2 => 
                           net75113, ZN => n48);
   U49 : AOI22_X1 port map( A1 => x(24), A2 => net75109, B1 => y(24), B2 => 
                           net75115, ZN => n49);
   U50 : AOI22_X1 port map( A1 => x(23), A2 => net75109, B1 => y(23), B2 => 
                           net75113, ZN => n50);
   U51 : AOI22_X1 port map( A1 => x(22), A2 => net75109, B1 => y(22), B2 => 
                           net75115, ZN => n51);
   U52 : AOI22_X1 port map( A1 => x(21), A2 => net75109, B1 => y(21), B2 => 
                           net75113, ZN => n52);
   U53 : AOI22_X1 port map( A1 => x(20), A2 => net75109, B1 => y(20), B2 => 
                           net75115, ZN => n53);
   U55 : AOI22_X1 port map( A1 => x(19), A2 => net75109, B1 => y(19), B2 => 
                           net75113, ZN => n55);
   U56 : AOI22_X1 port map( A1 => x(18), A2 => net75109, B1 => y(18), B2 => 
                           net75115, ZN => n56);
   U57 : AOI22_X1 port map( A1 => x(17), A2 => net75109, B1 => y(17), B2 => 
                           net75113, ZN => n57);
   U58 : AOI22_X1 port map( A1 => x(16), A2 => net75109, B1 => y(16), B2 => 
                           net75115, ZN => n58);
   U59 : AOI22_X1 port map( A1 => x(15), A2 => net75109, B1 => y(15), B2 => 
                           net75113, ZN => n59);
   U60 : AOI22_X1 port map( A1 => x(14), A2 => net75109, B1 => y(14), B2 => 
                           net75115, ZN => n60);
   U61 : AOI22_X1 port map( A1 => x(13), A2 => net75109, B1 => y(13), B2 => 
                           net75113, ZN => n61);
   U62 : AOI22_X1 port map( A1 => x(12), A2 => net75109, B1 => y(12), B2 => 
                           net75115, ZN => n62);
   U63 : AOI22_X1 port map( A1 => x(11), A2 => net75109, B1 => y(11), B2 => 
                           net75113, ZN => n63);
   U64 : AOI22_X1 port map( A1 => x(10), A2 => net75109, B1 => y(10), B2 => 
                           net75115, ZN => n64);
   U54 : AOI22_X1 port map( A1 => n68, A2 => x(1), B1 => n67, B2 => y(1), ZN =>
                           n54);
   U1 : NAND2_X1 port map( A1 => n68, A2 => x(0), ZN => n33);
   U2 : NAND2_X1 port map( A1 => n67, A2 => y(0), ZN => n65);
   U3 : NAND2_X1 port map( A1 => n65, A2 => n33, ZN => m(0));
   U5 : INV_X1 port map( A => sel, ZN => n68);
   U6 : INV_X1 port map( A => sel, ZN => net81028);
   U10 : INV_X1 port map( A => n40, ZN => m(3));
   U11 : INV_X2 port map( A => n39, ZN => m(4));
   U14 : INV_X1 port map( A => net81028, ZN => net82506);
   U17 : INV_X1 port map( A => n43, ZN => m(2));
   U22 : INV_X1 port map( A => n34, ZN => m(9));
   U23 : INV_X1 port map( A => n64, ZN => m(10));
   U24 : INV_X1 port map( A => n63, ZN => m(11));
   U25 : INV_X1 port map( A => n59, ZN => m(15));
   U26 : INV_X1 port map( A => n60, ZN => m(14));
   U27 : INV_X1 port map( A => n57, ZN => m(17));
   U28 : INV_X1 port map( A => n58, ZN => m(16));
   U29 : INV_X1 port map( A => n55, ZN => m(19));
   U30 : INV_X1 port map( A => n53, ZN => m(20));
   U31 : INV_X1 port map( A => n52, ZN => m(21));
   U32 : INV_X1 port map( A => n38, ZN => m(5));
   U33 : INV_X1 port map( A => n37, ZN => m(6));
   U65 : INV_X1 port map( A => n35, ZN => m(8));
   U66 : INV_X1 port map( A => n36, ZN => m(7));
   U67 : INV_X1 port map( A => n49, ZN => m(24));
   U68 : INV_X1 port map( A => n42, ZN => m(30));
   U69 : INV_X1 port map( A => n46, ZN => m(27));
   U70 : INV_X1 port map( A => n47, ZN => m(26));
   U71 : INV_X1 port map( A => n45, ZN => m(28));
   U72 : INV_X1 port map( A => n48, ZN => m(25));
   U73 : INV_X1 port map( A => n41, ZN => m(31));
   U74 : INV_X1 port map( A => n54, ZN => m(1));
   U4 : CLKBUF_X2 port map( A => net82506, Z => net75113);
   U7 : INV_X1 port map( A => net75113, ZN => net75109);
   U8 : BUF_X1 port map( A => net82506, Z => net75115);
   U9 : CLKBUF_X1 port map( A => n68, Z => net76536);
   U12 : BUF_X1 port map( A => sel, Z => n67);
   U13 : INV_X1 port map( A => n51, ZN => m(22));
   U15 : INV_X1 port map( A => n62, ZN => m(12));
   U16 : INV_X1 port map( A => n61, ZN => m(13));
   U18 : INV_X1 port map( A => n56, ZN => m(18));
   U19 : INV_X1 port map( A => n44, ZN => m(29));
   U20 : INV_X1 port map( A => n50, ZN => m(23));

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N1_0 is

   port( clk, rst, ld, data_in : in std_logic;  data_out : out std_logic);

end gen_reg_N1_0;

architecture SYN_behav of gen_reg_N1_0 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n3, B2 => ld, A => n2, ZN => n1);
   U3 : NAND2_X1 port map( A1 => ld, A2 => data_in, ZN => n2);
   data_out_reg_0_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           data_out, QN => n3);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity cond_branch is

   port( cond_in, jump_in, ctrl_in : in std_logic;  ctrl_out : out std_logic);

end cond_branch;

architecture SYN_dflow of cond_branch is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => ctrl_in, B => cond_in, ZN => n1);
   U1 : AND2_X1 port map( A1 => n1, A2 => jump_in, ZN => ctrl_out);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity zero_check_N32 is

   port( data_in : in std_logic_vector (31 downto 0);  ctrl_out : out std_logic
         );

end zero_check_N32;

architecture SYN_dflow of zero_check_N32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => 
                           ctrl_out);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => n4);
   U3 : NOR4_X1 port map( A1 => data_in(16), A2 => data_in(15), A3 => 
                           data_in(14), A4 => data_in(13), ZN => n6);
   U4 : NOR4_X1 port map( A1 => data_in(12), A2 => data_in(11), A3 => 
                           data_in(10), A4 => data_in(0), ZN => n5);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => n3);
   U6 : NOR4_X1 port map( A1 => data_in(23), A2 => data_in(22), A3 => 
                           data_in(21), A4 => data_in(20), ZN => n8);
   U7 : NOR4_X1 port map( A1 => data_in(1), A2 => data_in(19), A3 => 
                           data_in(18), A4 => data_in(17), ZN => n7);
   U8 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n2);
   U9 : NOR4_X1 port map( A1 => data_in(30), A2 => data_in(2), A3 => 
                           data_in(29), A4 => data_in(28), ZN => n10);
   U10 : NOR4_X1 port map( A1 => data_in(27), A2 => data_in(26), A3 => 
                           data_in(25), A4 => data_in(24), ZN => n9);
   U11 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n1);
   U12 : NOR4_X1 port map( A1 => data_in(9), A2 => data_in(8), A3 => data_in(7)
                           , A4 => data_in(6), ZN => n12);
   U13 : NOR4_X1 port map( A1 => data_in(5), A2 => data_in(4), A3 => data_in(3)
                           , A4 => data_in(31), ZN => n11);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_6 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_6;

architecture SYN_behav of gen_reg_N32_6 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n103, n104, n116, n117, n118, n119, n120, n121, n122, n123
      , n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n171, B2 => n103, A => n147, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n97, A2 => data_in(23), ZN => n147);
   U4 : OAI21_X1 port map( B1 => n172, B2 => n104, A => n146, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n97, ZN => n146);
   U6 : OAI21_X1 port map( B1 => n173, B2 => n103, A => n145, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => n104, ZN => n145);
   U8 : OAI21_X1 port map( B1 => n174, B2 => n103, A => n144, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => n104, ZN => n144);
   U10 : OAI21_X1 port map( B1 => n175, B2 => n103, A => n143, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => n97, ZN => n143);
   U12 : OAI21_X1 port map( B1 => n176, B2 => n104, A => n142, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => n97, ZN => n142);
   U14 : OAI21_X1 port map( B1 => n148, B2 => n104, A => n141, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => ld, ZN => n141);
   U16 : OAI21_X1 port map( B1 => n149, B2 => n104, A => n140, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n97, ZN => n140);
   U18 : OAI21_X1 port map( B1 => n150, B2 => n104, A => n139, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n97, ZN => n139);
   U20 : OAI21_X1 port map( B1 => n177, B2 => n103, A => n138, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n103, ZN => n138);
   U22 : OAI21_X1 port map( B1 => n151, B2 => n104, A => n137, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n97, ZN => n137);
   U24 : OAI21_X1 port map( B1 => n152, B2 => n104, A => n136, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n103, ZN => n136);
   U26 : OAI21_X1 port map( B1 => n153, B2 => n104, A => n135, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n97, ZN => n135);
   U28 : OAI21_X1 port map( B1 => n154, B2 => n103, A => n134, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => n97, ZN => n134);
   U30 : OAI21_X1 port map( B1 => n155, B2 => n97, A => n133, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => n97, ZN => n133);
   U32 : OAI21_X1 port map( B1 => n156, B2 => n103, A => n132, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n97, ZN => n132);
   U34 : OAI21_X1 port map( B1 => n157, B2 => n103, A => n131, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n103, ZN => n131);
   U36 : OAI21_X1 port map( B1 => n158, B2 => n103, A => n130, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n103, ZN => n130);
   U38 : OAI21_X1 port map( B1 => n159, B2 => n103, A => n129, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n97, ZN => n129);
   U40 : OAI21_X1 port map( B1 => n160, B2 => n104, A => n128, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => n97, ZN => n128);
   U42 : OAI21_X1 port map( B1 => n178, B2 => n104, A => n127, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => n97, ZN => n127);
   U44 : OAI21_X1 port map( B1 => n161, B2 => n104, A => n126, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => n97, ZN => n126);
   U46 : OAI21_X1 port map( B1 => n162, B2 => n103, A => n125, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => n103, ZN => n125);
   U48 : OAI21_X1 port map( B1 => n163, B2 => n103, A => n124, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => n97, ZN => n124);
   U50 : OAI21_X1 port map( B1 => n164, B2 => n104, A => n123, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n103, ZN => n123);
   U52 : OAI21_X1 port map( B1 => n165, B2 => n104, A => n122, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n97, ZN => n122);
   U54 : OAI21_X1 port map( B1 => n166, B2 => n103, A => n121, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n104, ZN => n121);
   U56 : OAI21_X1 port map( B1 => n167, B2 => n104, A => n120, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n97, ZN => n120);
   U58 : OAI21_X1 port map( B1 => n168, B2 => n103, A => n119, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n97, ZN => n119);
   U60 : OAI21_X1 port map( B1 => n169, B2 => n104, A => n118, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n97, ZN => n118);
   U62 : OAI21_X1 port map( B1 => n170, B2 => n103, A => n117, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => n104, ZN => n117);
   U64 : OAI21_X1 port map( B1 => n179, B2 => n104, A => n116, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n104, ZN => n116);
   U67 : CLKBUF_X1 port map( A => ld, Z => n97);
   U74 : CLKBUF_X1 port map( A => ld, Z => n103);
   U75 : CLKBUF_X1 port map( A => ld, Z => n104);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n179);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n178);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n177);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n176);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n175);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n174);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n173);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n172);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n171);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n170);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n169);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n168);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n167);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n166);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n165);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n164);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n163);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n162);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n161);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n160);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n159);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n158);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n157);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n156);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n155);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n154);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n153);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n152);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n151);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n150);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n149);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n148);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_mux21_N5 is

   port( sel : in std_logic;  x, y : in std_logic_vector (4 downto 0);  m : out
         std_logic_vector (4 downto 0));

end gen_mux21_N5;

architecture SYN_dflow of gen_mux21_N5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n16 : std_logic;

begin
   
   U7 : AOI22_X1 port map( A1 => x(4), A2 => n16, B1 => y(4), B2 => sel, ZN => 
                           n7);
   U8 : AOI22_X1 port map( A1 => x(3), A2 => n16, B1 => y(3), B2 => sel, ZN => 
                           n8);
   U9 : AOI22_X1 port map( A1 => x(2), A2 => n16, B1 => y(2), B2 => sel, ZN => 
                           n9);
   U10 : AOI22_X1 port map( A1 => x(1), A2 => n16, B1 => y(1), B2 => sel, ZN =>
                           n10);
   U11 : AOI22_X1 port map( A1 => x(0), A2 => n16, B1 => y(0), B2 => sel, ZN =>
                           n11);
   U1 : INV_X1 port map( A => n11, ZN => m(0));
   U2 : INV_X1 port map( A => sel, ZN => n16);
   U3 : INV_X1 port map( A => n10, ZN => m(1));
   U4 : INV_X1 port map( A => n9, ZN => m(2));
   U5 : INV_X1 port map( A => n8, ZN => m(3));
   U6 : INV_X1 port map( A => n7, ZN => m(4));

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity sign_ext_N_IN026_N_IN116_N_OUT32 is

   port( ctrl_in, zero_padding : in std_logic;  data_in : in std_logic_vector 
         (25 downto 0);  data_ext : out std_logic_vector (31 downto 0));

end sign_ext_N_IN026_N_IN116_N_OUT32;

architecture SYN_dflow of sign_ext_N_IN026_N_IN116_N_OUT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal data_ext_31_port, data_ext_24_port, data_ext_23_port, 
      data_ext_22_port, data_ext_21_port, data_ext_20_port, data_ext_19_port, 
      data_ext_18_port, data_ext_17_port, data_ext_16_port, n2, n3, n4, n5, n6,
      n7, n8, n9, n10, n11, n12, n13, n14 : std_logic;

begin
   data_ext <= ( data_ext_31_port, data_ext_31_port, data_ext_31_port, 
      data_ext_31_port, data_ext_31_port, data_ext_31_port, data_ext_31_port, 
      data_ext_24_port, data_ext_23_port, data_ext_22_port, data_ext_21_port, 
      data_ext_20_port, data_ext_19_port, data_ext_18_port, data_ext_17_port, 
      data_ext_16_port, data_in(15), data_in(14), data_in(13), data_in(12), 
      data_in(11), data_in(10), data_in(9), data_in(8), data_in(7), data_in(6),
      data_in(5), data_in(4), data_in(3), data_in(2), data_in(1), data_in(0) );
   
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => data_ext_31_port);
   U4 : NAND2_X1 port map( A1 => data_in(25), A2 => n14, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n2, A2 => n4, ZN => data_ext_24_port);
   U6 : NAND2_X1 port map( A1 => data_in(24), A2 => n14, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n5, ZN => data_ext_23_port);
   U8 : NAND2_X1 port map( A1 => data_in(23), A2 => n14, ZN => n5);
   U9 : NAND2_X1 port map( A1 => n2, A2 => n6, ZN => data_ext_22_port);
   U10 : NAND2_X1 port map( A1 => data_in(22), A2 => n14, ZN => n6);
   U11 : NAND2_X1 port map( A1 => n2, A2 => n7, ZN => data_ext_21_port);
   U12 : NAND2_X1 port map( A1 => data_in(21), A2 => n14, ZN => n7);
   U13 : NAND2_X1 port map( A1 => n2, A2 => n8, ZN => data_ext_20_port);
   U14 : NAND2_X1 port map( A1 => data_in(20), A2 => n14, ZN => n8);
   U15 : NAND2_X1 port map( A1 => n2, A2 => n9, ZN => data_ext_19_port);
   U16 : NAND2_X1 port map( A1 => data_in(19), A2 => n14, ZN => n9);
   U17 : NAND2_X1 port map( A1 => n2, A2 => n10, ZN => data_ext_18_port);
   U18 : NAND2_X1 port map( A1 => data_in(18), A2 => n14, ZN => n10);
   U19 : NAND2_X1 port map( A1 => n2, A2 => n11, ZN => data_ext_17_port);
   U20 : NAND2_X1 port map( A1 => data_in(17), A2 => n14, ZN => n11);
   U21 : NAND2_X1 port map( A1 => n2, A2 => n12, ZN => data_ext_16_port);
   U22 : NAND2_X1 port map( A1 => data_in(16), A2 => n14, ZN => n12);
   U23 : NAND2_X1 port map( A1 => n13, A2 => data_in(15), ZN => n2);
   U24 : NOR2_X1 port map( A1 => zero_padding, A2 => n14, ZN => n13);
   U2 : INV_X1 port map( A => ctrl_in, ZN => n14);

end SYN_dflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity reg_file_Dbits32_Abits5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end reg_file_Dbits32_Abits5;

architecture SYN_INTEGER of reg_file_Dbits32_Abits5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
      n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
      n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, 
      n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, 
      n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
      n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, 
      n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, 
      n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, 
      n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
      n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, 
      n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
      n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
      n3769, n3770, n3771, n3772, n3773, n3806, n3807, n3808, n3809, n3810, 
      n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, 
      n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, 
      n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, 
      n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, 
      n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
      n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3998, 
      n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
      n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
      n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
      n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
      n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, 
      n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
      n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
      n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n2130, n2135, n2140
      , n2145, n2150, n2155, n2160, n2165, n2170, n2175, n2180, n2185, n2190, 
      n2195, n2200, n2205, n2210, n2215, n2220, n2225, n2230, n2235, n2240, 
      n2245, n2250, n2255, n2260, n2265, n2270, n2352, n2355, n2358, n2361, 
      n2364, n2367, n2370, n2373, n2376, n2379, n2382, n2807, n2808, n2809, 
      n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
      n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
      n2830, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
      n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
      n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3802, n3803, n3804, n3805, n3870, n3871, n3872, n3873, n3874, n3875, 
      n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, 
      n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, 
      n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, 
      n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, 
      n3916, n3917, n3918, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1487, n1488, n1489, n1490, n1491, 
      n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
      n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
      n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, 
      n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, 
      n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, 
      n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, 
      n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, 
      n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
      n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, 
      n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, 
      n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, 
      n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, 
      n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, 
      n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, 
      n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, 
      n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, 
      n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, 
      n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, 
      n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, 
      n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, 
      n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
      n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, 
      n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, 
      n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
      n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
      n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, 
      n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
      n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
      n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, 
      n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, 
      n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, 
      n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, 
      n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, 
      n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, 
      n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, 
      n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, 
      n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, 
      n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
      n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, 
      n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, 
      n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, 
      n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, 
      n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, 
      n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, 
      n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
      n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, 
      n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, 
      n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, 
      n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, 
      n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, 
      n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, 
      n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, 
      n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, 
      n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, 
      n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, 
      n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, 
      n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, 
      n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2131, n2132, 
      n2133, n2134, n2136, n2137, n2138, n2139, n2141, n2142, n2143, n2144, 
      n2146, n2147, n2148, n2149, n2151, n2152, n2153, n2154, n2156, n2157, 
      n2158, n2159, n2161, n2162, n2163, n2164, n2166, n2167, n2168, n2169, 
      n2171, n2172, n2173, n2174, n2176, n2177, n2178, n2179, n2181, n2182, 
      n2183, n2184, n2186, n2187, n2188, n2189, n2191, n2192, n2193, n2194, 
      n2196, n2197, n2198, n2199, n2201, n2202, n2203, n2204, n2206, n2207, 
      n2208, n2209, n2211, n2212, n2213, n2214, n2216, n2217, n2218, n2219, 
      n2221, n2222, n2223, n2224, n2226, n2227, n2228, n2229, n2231, n2232, 
      n2233, n2234, n2236, n2237, n2238, n2239, n2241, n2242, n2243, n2244, 
      n2246, n2247, n2248, n2249, n2251, n2252, n2253, n2254, n2256, n2257, 
      n2258, n2259, n2261, n2262, n2263, n2264, n2266, n2267, n2268, n2269, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2353, n2354, n2356, n2357, n2359, n2360, n2362, n2363, n2365, 
      n2366, n2368, n2369, n2371, n2372, n2374, n2375, n2377, n2378, n2380, 
      n2381, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, 
      n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
      n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, 
      n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, 
      n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, 
      n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, 
      n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, 
      n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, 
      n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, 
      n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, 
      n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, 
      n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, 
      n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, 
      n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, 
      n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
      n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
      n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, 
      n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, 
      n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, 
      n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, 
      n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
      n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
      n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, 
      n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, 
      n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
      n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
      n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, 
      n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, 
      n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, 
      n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, 
      n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
      n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
      n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, 
      n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, 
      n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, 
      n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, 
      n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, 
      n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, 
      n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, 
      n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
      n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
      n2802, n2803, n2804, n2805, n2806, n2831, n2832, n2833, n2834, n2835, 
      n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, 
      n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, 
      n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, 
      n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, 
      n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
      n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, 
      n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, 
      n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
      n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, 
      n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, 
      n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, 
      n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, 
      n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, 
      n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
      n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, 
      n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, 
      n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
      n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
      n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
      n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, 
      n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3919, 
      n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, 
      n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
      n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
      n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
      n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
      n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, 
      n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, 
      n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n4190, n4191, 
      n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, 
      n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, 
      n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, 
      n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, 
      n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, 
      n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, 
      n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, 
      n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, 
      n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, 
      n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, 
      n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, 
      n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, 
      n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, 
      n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, 
      n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
      n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, 
      n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, 
      n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, 
      n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, 
      n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, 
      n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, 
      n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, 
      n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, 
      n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
      n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, 
      n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, 
      n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
      n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, 
      n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, 
      n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
      n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5335, 
      n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
      n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, 
      n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, 
      n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, 
      n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
      n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, 
      n5456, n5459, n5462, n5465, n5468, n5471, n5474, n5477, n5480, n5481, 
      n5486, n5489, n5492, n5495, n5498, n5499, n5504, n5506, n5509, n5513, 
      n5516, n5519, n5522, n5523, n5528, n5531, n5534, n5537, n5540, n5543, 
      n5546, n5549, n5552, n5556, n5557, n5562, n5564, n5565, n5567, n5573, 
      n5576, n5577, n5581, n5585, n5588, n5591, n5594, n5597, n5600, n5601, 
      n5605, n5609, n5612, n5615, n5618, n5621, n5624, n5627, n5629, n5633, 
      n5636, n5639, n5642, n5645, n5648, n5649, n5654, n5657, n5660, n5663, 
      n5666, n5669, n5672, n5673, n5677, n5681, n5684, n5687, n5690, n5693, 
      n5696, n5697, n5701, n5705, n5708, n5711, n5714, n5717, n5720, n5723, 
      n5725, n5729, n5732, n5735, n5738, n5741, n5744, n5745, n5750, n5753, 
      n5756, n5759, n5762, n5764, n5768, n5773, n5774, n5775, n5777, n5785, 
      n5786, n5790, n5791, n5793, n5795, n5803, n5804, n5808, n5809, n5812, 
      n5816, n5818, n5822, n5827, n5828, n5829, n5831, n5839, n5840, n5845, 
      n5846, n5850, n5851, n5854, n5858, n5863, n5864, n5868, n5869, n5871, 
      n5873, n5880, n5882, n5886, n5887, n5890, n5894, n5898, n5900, n5904, 
      n5906, n5907, n5909, n5916, n5918, n5922, n5923, n5925, n5930, n5932, 
      n5934, n5935, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, 
      n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, 
      n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, 
      n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, 
      n6085, n6086, n6087, n6088, n6089, n6090, n6603, n6604, n6605, n6606, 
      n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, 
      n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, 
      n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, 
      n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, 
      n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, 
      n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, 
      n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, 
      n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, 
      n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, 
      n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, 
      n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, 
      n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, 
      n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, 
      n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, 
      n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, 
      n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, 
      n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, 
      n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, 
      n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, 
      n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, 
      n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, 
      n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, 
      n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, 
      n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, 
      n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, 
      n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, 
      n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, 
      n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, 
      n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, 
      n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, 
      n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, 
      n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, 
      n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, 
      n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, 
      n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, 
      n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, 
      n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, 
      n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, 
      n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, 
      n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, 
      n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, 
      n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, 
      n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, 
      n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, 
      n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, 
      n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, 
      n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, 
      n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, 
      n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, 
      n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, 
      n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, 
      n7117, n7118, n7119, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, 
      n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, 
      n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, 
      n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, 
      n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, 
      n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, 
      n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, 
      n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, 
      n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, 
      n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, 
      n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, 
      n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, 
      n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, 
      n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, 
      n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, 
      n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, 
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, 
      n_2096 : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   U560 : OAI21_X1 port map( B1 => n5925, B2 => n5459, A => n1488, ZN => n4189)
                           ;
   U561 : NAND2_X1 port map( A1 => n5930, A2 => n7083, ZN => n1488);
   U562 : OAI21_X1 port map( B1 => n5925, B2 => n5462, A => n1489, ZN => n4188)
                           ;
   U563 : NAND2_X1 port map( A1 => n5930, A2 => n7082, ZN => n1489);
   U564 : OAI21_X1 port map( B1 => n5925, B2 => n5465, A => n1490, ZN => n4187)
                           ;
   U565 : NAND2_X1 port map( A1 => n5930, A2 => n7081, ZN => n1490);
   U566 : OAI21_X1 port map( B1 => n5925, B2 => n5468, A => n1491, ZN => n4186)
                           ;
   U567 : NAND2_X1 port map( A1 => n5925, A2 => n7080, ZN => n1491);
   U568 : OAI21_X1 port map( B1 => n5925, B2 => n5471, A => n1492, ZN => n4185)
                           ;
   U569 : NAND2_X1 port map( A1 => n5930, A2 => n7079, ZN => n1492);
   U570 : OAI21_X1 port map( B1 => n5925, B2 => n5474, A => n1493, ZN => n4184)
                           ;
   U571 : NAND2_X1 port map( A1 => n5925, A2 => n7078, ZN => n1493);
   U572 : OAI21_X1 port map( B1 => n5925, B2 => n5477, A => n1494, ZN => n4183)
                           ;
   U573 : NAND2_X1 port map( A1 => n5930, A2 => n7077, ZN => n1494);
   U574 : OAI21_X1 port map( B1 => n5925, B2 => n5480, A => n1495, ZN => n4182)
                           ;
   U575 : NAND2_X1 port map( A1 => n5925, A2 => n7076, ZN => n1495);
   U576 : OAI21_X1 port map( B1 => n5925, B2 => n6067, A => n1496, ZN => n4181)
                           ;
   U577 : NAND2_X1 port map( A1 => n5930, A2 => n7075, ZN => n1496);
   U578 : OAI21_X1 port map( B1 => n5925, B2 => n5486, A => n1497, ZN => n4180)
                           ;
   U579 : NAND2_X1 port map( A1 => n1487, A2 => n7074, ZN => n1497);
   U580 : OAI21_X1 port map( B1 => n5925, B2 => n5489, A => n1498, ZN => n4179)
                           ;
   U581 : NAND2_X1 port map( A1 => n5925, A2 => n7073, ZN => n1498);
   U582 : OAI21_X1 port map( B1 => n5925, B2 => n5492, A => n1499, ZN => n4178)
                           ;
   U583 : NAND2_X1 port map( A1 => n1487, A2 => n7072, ZN => n1499);
   U584 : OAI21_X1 port map( B1 => n5925, B2 => n5495, A => n1500, ZN => n4177)
                           ;
   U585 : NAND2_X1 port map( A1 => n1487, A2 => n7071, ZN => n1500);
   U586 : OAI21_X1 port map( B1 => n5930, B2 => n5498, A => n1501, ZN => n4176)
                           ;
   U587 : NAND2_X1 port map( A1 => n1487, A2 => n7070, ZN => n1501);
   U588 : OAI21_X1 port map( B1 => n5925, B2 => n6073, A => n1502, ZN => n4175)
                           ;
   U589 : NAND2_X1 port map( A1 => n1487, A2 => n7069, ZN => n1502);
   U590 : OAI21_X1 port map( B1 => n5930, B2 => n5504, A => n1503, ZN => n4174)
                           ;
   U591 : NAND2_X1 port map( A1 => n1487, A2 => n7068, ZN => n1503);
   U592 : OAI21_X1 port map( B1 => n5925, B2 => n6075, A => n1504, ZN => n4173)
                           ;
   U593 : NAND2_X1 port map( A1 => n1487, A2 => n7067, ZN => n1504);
   U594 : OAI21_X1 port map( B1 => n5930, B2 => n5509, A => n1505, ZN => n4172)
                           ;
   U595 : NAND2_X1 port map( A1 => n1487, A2 => n7066, ZN => n1505);
   U596 : OAI21_X1 port map( B1 => n5930, B2 => n5513, A => n1506, ZN => n4171)
                           ;
   U597 : NAND2_X1 port map( A1 => n5930, A2 => n7065, ZN => n1506);
   U598 : OAI21_X1 port map( B1 => n5930, B2 => n5516, A => n1507, ZN => n4170)
                           ;
   U599 : NAND2_X1 port map( A1 => n1487, A2 => n7064, ZN => n1507);
   U600 : OAI21_X1 port map( B1 => n5930, B2 => n5519, A => n1508, ZN => n4169)
                           ;
   U601 : NAND2_X1 port map( A1 => n1487, A2 => n7063, ZN => n1508);
   U602 : OAI21_X1 port map( B1 => n5930, B2 => n5522, A => n1509, ZN => n4168)
                           ;
   U603 : NAND2_X1 port map( A1 => n5930, A2 => n7062, ZN => n1509);
   U604 : OAI21_X1 port map( B1 => n5930, B2 => n6081, A => n1510, ZN => n4167)
                           ;
   U605 : NAND2_X1 port map( A1 => n1487, A2 => n7061, ZN => n1510);
   U606 : OAI21_X1 port map( B1 => n1487, B2 => n5528, A => n1511, ZN => n4166)
                           ;
   U607 : NAND2_X1 port map( A1 => n1487, A2 => n7060, ZN => n1511);
   U608 : OAI21_X1 port map( B1 => n5930, B2 => n5531, A => n1512, ZN => n4165)
                           ;
   U609 : NAND2_X1 port map( A1 => n1487, A2 => n7059, ZN => n1512);
   U610 : OAI21_X1 port map( B1 => n1487, B2 => n5534, A => n1513, ZN => n4164)
                           ;
   U611 : NAND2_X1 port map( A1 => n1487, A2 => n7058, ZN => n1513);
   U612 : OAI21_X1 port map( B1 => n1487, B2 => n5537, A => n1514, ZN => n4163)
                           ;
   U613 : NAND2_X1 port map( A1 => n1487, A2 => n7057, ZN => n1514);
   U614 : OAI21_X1 port map( B1 => n1487, B2 => n5540, A => n1515, ZN => n4162)
                           ;
   U615 : NAND2_X1 port map( A1 => n1487, A2 => n7056, ZN => n1515);
   U616 : OAI21_X1 port map( B1 => n1487, B2 => n5543, A => n1516, ZN => n4161)
                           ;
   U617 : NAND2_X1 port map( A1 => n1487, A2 => n7055, ZN => n1516);
   U618 : OAI21_X1 port map( B1 => n1487, B2 => n5546, A => n1517, ZN => n4160)
                           ;
   U619 : NAND2_X1 port map( A1 => n1487, A2 => n7054, ZN => n1517);
   U620 : OAI21_X1 port map( B1 => n5930, B2 => n5549, A => n1518, ZN => n4159)
                           ;
   U621 : NAND2_X1 port map( A1 => n5930, A2 => n7053, ZN => n1518);
   U622 : OAI21_X1 port map( B1 => n5925, B2 => n5552, A => n1519, ZN => n4158)
                           ;
   U623 : NAND2_X1 port map( A1 => n5930, A2 => n7052, ZN => n1519);
   U624 : NAND2_X1 port map( A1 => n1520, A2 => n1521, ZN => n1487);
   U625 : OAI21_X1 port map( B1 => n5459, B2 => n5922, A => n1523, ZN => n4157)
                           ;
   U626 : NAND2_X1 port map( A1 => n5923, A2 => n6710, ZN => n1523);
   U627 : OAI21_X1 port map( B1 => n5462, B2 => n5923, A => n1524, ZN => n4156)
                           ;
   U628 : NAND2_X1 port map( A1 => n5923, A2 => n6709, ZN => n1524);
   U629 : OAI21_X1 port map( B1 => n5465, B2 => n5922, A => n1525, ZN => n4155)
                           ;
   U630 : NAND2_X1 port map( A1 => n5922, A2 => n6708, ZN => n1525);
   U631 : OAI21_X1 port map( B1 => n5468, B2 => n5922, A => n1526, ZN => n4154)
                           ;
   U632 : NAND2_X1 port map( A1 => n2270, A2 => n1522, ZN => n1526);
   U633 : OAI21_X1 port map( B1 => n5471, B2 => n5923, A => n1527, ZN => n4153)
                           ;
   U634 : NAND2_X1 port map( A1 => n2265, A2 => n5922, ZN => n1527);
   U635 : OAI21_X1 port map( B1 => n5474, B2 => n5922, A => n1528, ZN => n4152)
                           ;
   U636 : NAND2_X1 port map( A1 => n2260, A2 => n1522, ZN => n1528);
   U637 : OAI21_X1 port map( B1 => n5477, B2 => n5922, A => n1529, ZN => n4151)
                           ;
   U638 : NAND2_X1 port map( A1 => n2255, A2 => n1522, ZN => n1529);
   U639 : OAI21_X1 port map( B1 => n5480, B2 => n5922, A => n1530, ZN => n4150)
                           ;
   U640 : NAND2_X1 port map( A1 => n2250, A2 => n1522, ZN => n1530);
   U641 : OAI21_X1 port map( B1 => n6067, B2 => n5922, A => n1531, ZN => n4149)
                           ;
   U642 : NAND2_X1 port map( A1 => n2245, A2 => n5922, ZN => n1531);
   U643 : OAI21_X1 port map( B1 => n5486, B2 => n5922, A => n1532, ZN => n4148)
                           ;
   U644 : NAND2_X1 port map( A1 => n2240, A2 => n1522, ZN => n1532);
   U645 : OAI21_X1 port map( B1 => n5489, B2 => n5922, A => n1533, ZN => n4147)
                           ;
   U646 : NAND2_X1 port map( A1 => n2235, A2 => n1522, ZN => n1533);
   U647 : OAI21_X1 port map( B1 => n5492, B2 => n5922, A => n1534, ZN => n4146)
                           ;
   U648 : NAND2_X1 port map( A1 => n2230, A2 => n5923, ZN => n1534);
   U649 : OAI21_X1 port map( B1 => n5495, B2 => n5922, A => n1535, ZN => n4145)
                           ;
   U650 : NAND2_X1 port map( A1 => n2225, A2 => n5922, ZN => n1535);
   U651 : OAI21_X1 port map( B1 => n5498, B2 => n5922, A => n1536, ZN => n4144)
                           ;
   U652 : NAND2_X1 port map( A1 => n2220, A2 => n1522, ZN => n1536);
   U653 : OAI21_X1 port map( B1 => n6073, B2 => n5922, A => n1537, ZN => n4143)
                           ;
   U654 : NAND2_X1 port map( A1 => n2215, A2 => n5923, ZN => n1537);
   U655 : OAI21_X1 port map( B1 => n5504, B2 => n5923, A => n1538, ZN => n4142)
                           ;
   U656 : NAND2_X1 port map( A1 => n2210, A2 => n5923, ZN => n1538);
   U657 : OAI21_X1 port map( B1 => n6075, B2 => n5923, A => n1539, ZN => n4141)
                           ;
   U658 : NAND2_X1 port map( A1 => n2205, A2 => n1522, ZN => n1539);
   U659 : OAI21_X1 port map( B1 => n5509, B2 => n5923, A => n1540, ZN => n4140)
                           ;
   U660 : NAND2_X1 port map( A1 => n2200, A2 => n1522, ZN => n1540);
   U661 : OAI21_X1 port map( B1 => n5513, B2 => n5923, A => n1541, ZN => n4139)
                           ;
   U662 : NAND2_X1 port map( A1 => n2195, A2 => n1522, ZN => n1541);
   U663 : OAI21_X1 port map( B1 => n5516, B2 => n5923, A => n1542, ZN => n4138)
                           ;
   U664 : NAND2_X1 port map( A1 => n2190, A2 => n1522, ZN => n1542);
   U665 : OAI21_X1 port map( B1 => n5519, B2 => n5923, A => n1543, ZN => n4137)
                           ;
   U666 : NAND2_X1 port map( A1 => n2185, A2 => n1522, ZN => n1543);
   U667 : OAI21_X1 port map( B1 => n5522, B2 => n5923, A => n1544, ZN => n4136)
                           ;
   U668 : NAND2_X1 port map( A1 => n2180, A2 => n1522, ZN => n1544);
   U669 : OAI21_X1 port map( B1 => n6081, B2 => n5923, A => n1545, ZN => n4135)
                           ;
   U670 : NAND2_X1 port map( A1 => n2175, A2 => n1522, ZN => n1545);
   U671 : OAI21_X1 port map( B1 => n5528, B2 => n5923, A => n1546, ZN => n4134)
                           ;
   U672 : NAND2_X1 port map( A1 => n2170, A2 => n1522, ZN => n1546);
   U673 : OAI21_X1 port map( B1 => n5531, B2 => n5923, A => n1547, ZN => n4133)
                           ;
   U674 : NAND2_X1 port map( A1 => n2165, A2 => n1522, ZN => n1547);
   U675 : OAI21_X1 port map( B1 => n5534, B2 => n5923, A => n1548, ZN => n4132)
                           ;
   U676 : NAND2_X1 port map( A1 => n2160, A2 => n1522, ZN => n1548);
   U677 : OAI21_X1 port map( B1 => n5537, B2 => n5923, A => n1549, ZN => n4131)
                           ;
   U678 : NAND2_X1 port map( A1 => n2155, A2 => n1522, ZN => n1549);
   U679 : OAI21_X1 port map( B1 => n5540, B2 => n5923, A => n1550, ZN => n4130)
                           ;
   U680 : NAND2_X1 port map( A1 => n2150, A2 => n1522, ZN => n1550);
   U681 : OAI21_X1 port map( B1 => n5543, B2 => n5922, A => n1551, ZN => n4129)
                           ;
   U682 : NAND2_X1 port map( A1 => n2145, A2 => n1522, ZN => n1551);
   U683 : OAI21_X1 port map( B1 => n5546, B2 => n5923, A => n1552, ZN => n4128)
                           ;
   U684 : NAND2_X1 port map( A1 => n2140, A2 => n1522, ZN => n1552);
   U685 : OAI21_X1 port map( B1 => n5549, B2 => n5922, A => n1553, ZN => n4127)
                           ;
   U686 : NAND2_X1 port map( A1 => n2135, A2 => n1522, ZN => n1553);
   U687 : OAI21_X1 port map( B1 => n5552, B2 => n5922, A => n1554, ZN => n4126)
                           ;
   U688 : NAND2_X1 port map( A1 => n2130, A2 => n1522, ZN => n1554);
   U689 : NAND2_X1 port map( A1 => n1555, A2 => n1556, ZN => n1522);
   U690 : OAI21_X1 port map( B1 => n5459, B2 => n5916, A => n1558, ZN => n4125)
                           ;
   U691 : NAND2_X1 port map( A1 => n1557, A2 => n7051, ZN => n1558);
   U692 : OAI21_X1 port map( B1 => n5462, B2 => n1557, A => n1559, ZN => n4124)
                           ;
   U693 : NAND2_X1 port map( A1 => n1557, A2 => n7050, ZN => n1559);
   U694 : OAI21_X1 port map( B1 => n5465, B2 => n5916, A => n1560, ZN => n4123)
                           ;
   U695 : NAND2_X1 port map( A1 => n1557, A2 => n7049, ZN => n1560);
   U696 : OAI21_X1 port map( B1 => n5468, B2 => n1557, A => n1561, ZN => n4122)
                           ;
   U697 : NAND2_X1 port map( A1 => n1557, A2 => n7048, ZN => n1561);
   U698 : OAI21_X1 port map( B1 => n5471, B2 => n1557, A => n1562, ZN => n4121)
                           ;
   U699 : NAND2_X1 port map( A1 => n5918, A2 => n7047, ZN => n1562);
   U700 : OAI21_X1 port map( B1 => n5474, B2 => n5916, A => n1563, ZN => n4120)
                           ;
   U701 : NAND2_X1 port map( A1 => n1557, A2 => n7046, ZN => n1563);
   U702 : OAI21_X1 port map( B1 => n5477, B2 => n5916, A => n1564, ZN => n4119)
                           ;
   U703 : NAND2_X1 port map( A1 => n1557, A2 => n7045, ZN => n1564);
   U704 : OAI21_X1 port map( B1 => n5480, B2 => n5916, A => n1565, ZN => n4118)
                           ;
   U705 : NAND2_X1 port map( A1 => n1557, A2 => n7044, ZN => n1565);
   U706 : OAI21_X1 port map( B1 => n6067, B2 => n5916, A => n1566, ZN => n4117)
                           ;
   U707 : NAND2_X1 port map( A1 => n1557, A2 => n7043, ZN => n1566);
   U708 : OAI21_X1 port map( B1 => n5486, B2 => n5916, A => n1567, ZN => n4116)
                           ;
   U709 : NAND2_X1 port map( A1 => n1557, A2 => n7042, ZN => n1567);
   U710 : OAI21_X1 port map( B1 => n5489, B2 => n5916, A => n1568, ZN => n4115)
                           ;
   U711 : NAND2_X1 port map( A1 => n1557, A2 => n7041, ZN => n1568);
   U712 : OAI21_X1 port map( B1 => n5492, B2 => n5916, A => n1569, ZN => n4114)
                           ;
   U713 : NAND2_X1 port map( A1 => n1557, A2 => n7040, ZN => n1569);
   U714 : OAI21_X1 port map( B1 => n5495, B2 => n5916, A => n1570, ZN => n4113)
                           ;
   U715 : NAND2_X1 port map( A1 => n1557, A2 => n7039, ZN => n1570);
   U716 : OAI21_X1 port map( B1 => n5498, B2 => n5916, A => n1571, ZN => n4112)
                           ;
   U717 : NAND2_X1 port map( A1 => n1557, A2 => n7038, ZN => n1571);
   U718 : OAI21_X1 port map( B1 => n6073, B2 => n5916, A => n1572, ZN => n4111)
                           ;
   U719 : NAND2_X1 port map( A1 => n5916, A2 => n7037, ZN => n1572);
   U720 : OAI21_X1 port map( B1 => n5504, B2 => n5918, A => n1573, ZN => n4110)
                           ;
   U721 : NAND2_X1 port map( A1 => n5916, A2 => n7036, ZN => n1573);
   U722 : OAI21_X1 port map( B1 => n6075, B2 => n5916, A => n1574, ZN => n4109)
                           ;
   U723 : NAND2_X1 port map( A1 => n5916, A2 => n7035, ZN => n1574);
   U724 : OAI21_X1 port map( B1 => n5509, B2 => n5918, A => n1575, ZN => n4108)
                           ;
   U725 : NAND2_X1 port map( A1 => n5918, A2 => n7034, ZN => n1575);
   U726 : OAI21_X1 port map( B1 => n5513, B2 => n5916, A => n1576, ZN => n4107)
                           ;
   U727 : NAND2_X1 port map( A1 => n5918, A2 => n7033, ZN => n1576);
   U728 : OAI21_X1 port map( B1 => n5516, B2 => n5918, A => n1577, ZN => n4106)
                           ;
   U729 : NAND2_X1 port map( A1 => n5918, A2 => n7032, ZN => n1577);
   U730 : OAI21_X1 port map( B1 => n5519, B2 => n5916, A => n1578, ZN => n4105)
                           ;
   U731 : NAND2_X1 port map( A1 => n5918, A2 => n7031, ZN => n1578);
   U732 : OAI21_X1 port map( B1 => n5522, B2 => n5918, A => n1579, ZN => n4104)
                           ;
   U733 : NAND2_X1 port map( A1 => n5918, A2 => n7030, ZN => n1579);
   U734 : OAI21_X1 port map( B1 => n6081, B2 => n5916, A => n1580, ZN => n4103)
                           ;
   U735 : NAND2_X1 port map( A1 => n5918, A2 => n7029, ZN => n1580);
   U736 : OAI21_X1 port map( B1 => n5528, B2 => n5918, A => n1581, ZN => n4102)
                           ;
   U737 : NAND2_X1 port map( A1 => n5918, A2 => n7028, ZN => n1581);
   U738 : OAI21_X1 port map( B1 => n5531, B2 => n5916, A => n1582, ZN => n4101)
                           ;
   U739 : NAND2_X1 port map( A1 => n5918, A2 => n7027, ZN => n1582);
   U740 : OAI21_X1 port map( B1 => n5534, B2 => n5918, A => n1583, ZN => n4100)
                           ;
   U741 : NAND2_X1 port map( A1 => n1557, A2 => n7026, ZN => n1583);
   U742 : OAI21_X1 port map( B1 => n5537, B2 => n1557, A => n1584, ZN => n4099)
                           ;
   U743 : NAND2_X1 port map( A1 => n5918, A2 => n7025, ZN => n1584);
   U744 : OAI21_X1 port map( B1 => n5540, B2 => n5918, A => n1585, ZN => n4098)
                           ;
   U745 : NAND2_X1 port map( A1 => n1557, A2 => n7024, ZN => n1585);
   U746 : OAI21_X1 port map( B1 => n5543, B2 => n5918, A => n1586, ZN => n4097)
                           ;
   U747 : NAND2_X1 port map( A1 => n1557, A2 => n7023, ZN => n1586);
   U748 : OAI21_X1 port map( B1 => n5546, B2 => n5918, A => n1587, ZN => n4096)
                           ;
   U749 : NAND2_X1 port map( A1 => n1557, A2 => n7022, ZN => n1587);
   U750 : OAI21_X1 port map( B1 => n5549, B2 => n5918, A => n1588, ZN => n4095)
                           ;
   U751 : NAND2_X1 port map( A1 => n1557, A2 => n7021, ZN => n1588);
   U752 : OAI21_X1 port map( B1 => n5552, B2 => n1557, A => n1589, ZN => n4094)
                           ;
   U753 : NAND2_X1 port map( A1 => n1557, A2 => n7020, ZN => n1589);
   U754 : NAND2_X1 port map( A1 => n1590, A2 => n1556, ZN => n1557);
   U755 : OAI21_X1 port map( B1 => n5459, B2 => n1591, A => n1592, ZN => n4093)
                           ;
   U756 : NAND2_X1 port map( A1 => n5907, A2 => n7019, ZN => n1592);
   U757 : OAI21_X1 port map( B1 => n5462, B2 => n5909, A => n1593, ZN => n4092)
                           ;
   U758 : NAND2_X1 port map( A1 => n5907, A2 => n7018, ZN => n1593);
   U759 : OAI21_X1 port map( B1 => n5465, B2 => n1591, A => n1594, ZN => n4091)
                           ;
   U760 : NAND2_X1 port map( A1 => n5907, A2 => n7017, ZN => n1594);
   U761 : OAI21_X1 port map( B1 => n5468, B2 => n5909, A => n1595, ZN => n4090)
                           ;
   U762 : NAND2_X1 port map( A1 => n5907, A2 => n7016, ZN => n1595);
   U763 : OAI21_X1 port map( B1 => n5471, B2 => n5909, A => n1596, ZN => n4089)
                           ;
   U764 : NAND2_X1 port map( A1 => n5907, A2 => n7015, ZN => n1596);
   U765 : OAI21_X1 port map( B1 => n5474, B2 => n1591, A => n1597, ZN => n4088)
                           ;
   U766 : NAND2_X1 port map( A1 => n5907, A2 => n7014, ZN => n1597);
   U767 : OAI21_X1 port map( B1 => n5477, B2 => n1591, A => n1598, ZN => n4087)
                           ;
   U768 : NAND2_X1 port map( A1 => n5909, A2 => n7013, ZN => n1598);
   U769 : OAI21_X1 port map( B1 => n5480, B2 => n1591, A => n1599, ZN => n4086)
                           ;
   U770 : NAND2_X1 port map( A1 => n5909, A2 => n7012, ZN => n1599);
   U771 : OAI21_X1 port map( B1 => n6067, B2 => n1591, A => n1600, ZN => n4085)
                           ;
   U772 : NAND2_X1 port map( A1 => n5909, A2 => n7011, ZN => n1600);
   U773 : OAI21_X1 port map( B1 => n5486, B2 => n1591, A => n1601, ZN => n4084)
                           ;
   U774 : NAND2_X1 port map( A1 => n5909, A2 => n7010, ZN => n1601);
   U775 : OAI21_X1 port map( B1 => n5489, B2 => n1591, A => n1602, ZN => n4083)
                           ;
   U776 : NAND2_X1 port map( A1 => n5909, A2 => n7009, ZN => n1602);
   U777 : OAI21_X1 port map( B1 => n5492, B2 => n1591, A => n1603, ZN => n4082)
                           ;
   U778 : NAND2_X1 port map( A1 => n5909, A2 => n7008, ZN => n1603);
   U779 : OAI21_X1 port map( B1 => n5495, B2 => n1591, A => n1604, ZN => n4081)
                           ;
   U780 : NAND2_X1 port map( A1 => n5909, A2 => n7007, ZN => n1604);
   U781 : OAI21_X1 port map( B1 => n5498, B2 => n1591, A => n1605, ZN => n4080)
                           ;
   U782 : NAND2_X1 port map( A1 => n5907, A2 => n7006, ZN => n1605);
   U783 : OAI21_X1 port map( B1 => n6073, B2 => n1591, A => n1606, ZN => n4079)
                           ;
   U784 : NAND2_X1 port map( A1 => n5909, A2 => n7005, ZN => n1606);
   U785 : OAI21_X1 port map( B1 => n5504, B2 => n5909, A => n1607, ZN => n4078)
                           ;
   U786 : NAND2_X1 port map( A1 => n5909, A2 => n7004, ZN => n1607);
   U787 : OAI21_X1 port map( B1 => n6075, B2 => n1591, A => n1608, ZN => n4077)
                           ;
   U788 : NAND2_X1 port map( A1 => n5909, A2 => n7003, ZN => n1608);
   U789 : OAI21_X1 port map( B1 => n5509, B2 => n5909, A => n1609, ZN => n4076)
                           ;
   U790 : NAND2_X1 port map( A1 => n5907, A2 => n7002, ZN => n1609);
   U791 : OAI21_X1 port map( B1 => n5513, B2 => n1591, A => n1610, ZN => n4075)
                           ;
   U792 : NAND2_X1 port map( A1 => n5909, A2 => n7001, ZN => n1610);
   U793 : OAI21_X1 port map( B1 => n5516, B2 => n5907, A => n1611, ZN => n4074)
                           ;
   U794 : NAND2_X1 port map( A1 => n5907, A2 => n7000, ZN => n1611);
   U795 : OAI21_X1 port map( B1 => n5519, B2 => n5909, A => n1612, ZN => n4073)
                           ;
   U796 : NAND2_X1 port map( A1 => n5909, A2 => n6999, ZN => n1612);
   U797 : OAI21_X1 port map( B1 => n5522, B2 => n1591, A => n1613, ZN => n4072)
                           ;
   U798 : NAND2_X1 port map( A1 => n5907, A2 => n6998, ZN => n1613);
   U799 : OAI21_X1 port map( B1 => n6081, B2 => n1591, A => n1614, ZN => n4071)
                           ;
   U800 : NAND2_X1 port map( A1 => n5909, A2 => n6997, ZN => n1614);
   U801 : OAI21_X1 port map( B1 => n5528, B2 => n1591, A => n1615, ZN => n4070)
                           ;
   U802 : NAND2_X1 port map( A1 => n5907, A2 => n6996, ZN => n1615);
   U803 : OAI21_X1 port map( B1 => n5531, B2 => n1591, A => n1616, ZN => n4069)
                           ;
   U804 : NAND2_X1 port map( A1 => n5907, A2 => n6995, ZN => n1616);
   U805 : OAI21_X1 port map( B1 => n5534, B2 => n1591, A => n1617, ZN => n4068)
                           ;
   U806 : NAND2_X1 port map( A1 => n5907, A2 => n6994, ZN => n1617);
   U807 : OAI21_X1 port map( B1 => n5537, B2 => n1591, A => n1618, ZN => n4067)
                           ;
   U808 : NAND2_X1 port map( A1 => n5907, A2 => n6993, ZN => n1618);
   U809 : OAI21_X1 port map( B1 => n5540, B2 => n1591, A => n1619, ZN => n4066)
                           ;
   U810 : NAND2_X1 port map( A1 => n5907, A2 => n6992, ZN => n1619);
   U811 : OAI21_X1 port map( B1 => n5543, B2 => n1591, A => n1620, ZN => n4065)
                           ;
   U812 : NAND2_X1 port map( A1 => n5907, A2 => n6991, ZN => n1620);
   U813 : OAI21_X1 port map( B1 => n5546, B2 => n1591, A => n1621, ZN => n4064)
                           ;
   U814 : NAND2_X1 port map( A1 => n5907, A2 => n6990, ZN => n1621);
   U815 : OAI21_X1 port map( B1 => n5549, B2 => n1591, A => n1622, ZN => n4063)
                           ;
   U816 : NAND2_X1 port map( A1 => n5907, A2 => n6989, ZN => n1622);
   U817 : OAI21_X1 port map( B1 => n5552, B2 => n5909, A => n1623, ZN => n4062)
                           ;
   U818 : NAND2_X1 port map( A1 => n5907, A2 => n6988, ZN => n1623);
   U819 : NAND2_X1 port map( A1 => n1624, A2 => n1556, ZN => n1591);
   U820 : OAI21_X1 port map( B1 => n5459, B2 => n5904, A => n1626, ZN => n4061)
                           ;
   U821 : NAND2_X1 port map( A1 => n2382, A2 => n1625, ZN => n1626);
   U822 : OAI21_X1 port map( B1 => n5462, B2 => n5906, A => n1627, ZN => n4060)
                           ;
   U823 : NAND2_X1 port map( A1 => n2379, A2 => n5906, ZN => n1627);
   U824 : OAI21_X1 port map( B1 => n5465, B2 => n5904, A => n1628, ZN => n4059)
                           ;
   U825 : NAND2_X1 port map( A1 => n2376, A2 => n1625, ZN => n1628);
   U826 : OAI21_X1 port map( B1 => n5468, B2 => n5904, A => n1629, ZN => n4058)
                           ;
   U827 : NAND2_X1 port map( A1 => n2373, A2 => n5906, ZN => n1629);
   U828 : OAI21_X1 port map( B1 => n5471, B2 => n5906, A => n1630, ZN => n4057)
                           ;
   U829 : NAND2_X1 port map( A1 => n2370, A2 => n5906, ZN => n1630);
   U830 : OAI21_X1 port map( B1 => n5474, B2 => n5904, A => n1631, ZN => n4056)
                           ;
   U831 : NAND2_X1 port map( A1 => n2367, A2 => n1625, ZN => n1631);
   U832 : OAI21_X1 port map( B1 => n5477, B2 => n5904, A => n1632, ZN => n4055)
                           ;
   U833 : NAND2_X1 port map( A1 => n2364, A2 => n5906, ZN => n1632);
   U834 : OAI21_X1 port map( B1 => n5480, B2 => n5904, A => n1633, ZN => n4054)
                           ;
   U835 : NAND2_X1 port map( A1 => n2361, A2 => n5906, ZN => n1633);
   U836 : OAI21_X1 port map( B1 => n6067, B2 => n5904, A => n1634, ZN => n4053)
                           ;
   U837 : NAND2_X1 port map( A1 => n2358, A2 => n5906, ZN => n1634);
   U838 : OAI21_X1 port map( B1 => n5486, B2 => n5904, A => n1635, ZN => n4052)
                           ;
   U839 : NAND2_X1 port map( A1 => n2355, A2 => n5906, ZN => n1635);
   U840 : OAI21_X1 port map( B1 => n5489, B2 => n5904, A => n1636, ZN => n4051)
                           ;
   U841 : NAND2_X1 port map( A1 => n2352, A2 => n5906, ZN => n1636);
   U842 : OAI21_X1 port map( B1 => n5492, B2 => n5904, A => n1637, ZN => n4050)
                           ;
   U843 : NAND2_X1 port map( A1 => n1625, A2 => n6763, ZN => n1637);
   U844 : OAI21_X1 port map( B1 => n5495, B2 => n5904, A => n1638, ZN => n4049)
                           ;
   U845 : NAND2_X1 port map( A1 => n1625, A2 => n6762, ZN => n1638);
   U846 : OAI21_X1 port map( B1 => n5498, B2 => n5904, A => n1639, ZN => n4048)
                           ;
   U847 : NAND2_X1 port map( A1 => n1625, A2 => n6761, ZN => n1639);
   U848 : OAI21_X1 port map( B1 => n6073, B2 => n5904, A => n1640, ZN => n4047)
                           ;
   U849 : NAND2_X1 port map( A1 => n1625, A2 => n6760, ZN => n1640);
   U850 : OAI21_X1 port map( B1 => n5504, B2 => n5904, A => n1641, ZN => n4046)
                           ;
   U851 : NAND2_X1 port map( A1 => n1625, A2 => n6759, ZN => n1641);
   U852 : OAI21_X1 port map( B1 => n6075, B2 => n5906, A => n1642, ZN => n4045)
                           ;
   U853 : NAND2_X1 port map( A1 => n1625, A2 => n6758, ZN => n1642);
   U854 : OAI21_X1 port map( B1 => n5509, B2 => n5904, A => n1643, ZN => n4044)
                           ;
   U855 : NAND2_X1 port map( A1 => n1625, A2 => n6757, ZN => n1643);
   U856 : OAI21_X1 port map( B1 => n5513, B2 => n5906, A => n1644, ZN => n4043)
                           ;
   U857 : NAND2_X1 port map( A1 => n1625, A2 => n6756, ZN => n1644);
   U858 : OAI21_X1 port map( B1 => n5516, B2 => n5904, A => n1645, ZN => n4042)
                           ;
   U859 : NAND2_X1 port map( A1 => n1625, A2 => n6755, ZN => n1645);
   U860 : OAI21_X1 port map( B1 => n5519, B2 => n5906, A => n1646, ZN => n4041)
                           ;
   U861 : NAND2_X1 port map( A1 => n1625, A2 => n6754, ZN => n1646);
   U862 : OAI21_X1 port map( B1 => n5522, B2 => n5904, A => n1647, ZN => n4040)
                           ;
   U863 : NAND2_X1 port map( A1 => n1625, A2 => n6753, ZN => n1647);
   U864 : OAI21_X1 port map( B1 => n6081, B2 => n5906, A => n1648, ZN => n4039)
                           ;
   U865 : NAND2_X1 port map( A1 => n1625, A2 => n6752, ZN => n1648);
   U866 : OAI21_X1 port map( B1 => n5528, B2 => n5904, A => n1649, ZN => n4038)
                           ;
   U867 : NAND2_X1 port map( A1 => n1625, A2 => n6751, ZN => n1649);
   U868 : OAI21_X1 port map( B1 => n5531, B2 => n5906, A => n1650, ZN => n4037)
                           ;
   U869 : NAND2_X1 port map( A1 => n1625, A2 => n6750, ZN => n1650);
   U870 : OAI21_X1 port map( B1 => n5534, B2 => n5904, A => n1651, ZN => n4036)
                           ;
   U871 : NAND2_X1 port map( A1 => n1625, A2 => n6749, ZN => n1651);
   U872 : OAI21_X1 port map( B1 => n5537, B2 => n5906, A => n1652, ZN => n4035)
                           ;
   U873 : NAND2_X1 port map( A1 => n1625, A2 => n6748, ZN => n1652);
   U874 : OAI21_X1 port map( B1 => n5540, B2 => n5906, A => n1653, ZN => n4034)
                           ;
   U875 : NAND2_X1 port map( A1 => n1625, A2 => n6747, ZN => n1653);
   U876 : OAI21_X1 port map( B1 => n5543, B2 => n5906, A => n1654, ZN => n4033)
                           ;
   U877 : NAND2_X1 port map( A1 => n5904, A2 => n6746, ZN => n1654);
   U878 : OAI21_X1 port map( B1 => n5546, B2 => n5906, A => n1655, ZN => n4032)
                           ;
   U879 : NAND2_X1 port map( A1 => n1625, A2 => n6745, ZN => n1655);
   U880 : OAI21_X1 port map( B1 => n5549, B2 => n5906, A => n1656, ZN => n4031)
                           ;
   U881 : NAND2_X1 port map( A1 => n1625, A2 => n6744, ZN => n1656);
   U882 : OAI21_X1 port map( B1 => n5552, B2 => n1625, A => n1657, ZN => n4030)
                           ;
   U883 : NAND2_X1 port map( A1 => n1625, A2 => n6743, ZN => n1657);
   U884 : NAND2_X1 port map( A1 => n1658, A2 => n1556, ZN => n1625);
   U885 : OAI21_X1 port map( B1 => n5459, B2 => n5898, A => n1660, ZN => n4029)
                           ;
   U886 : NAND2_X1 port map( A1 => n1659, A2 => n6707, ZN => n1660);
   U887 : OAI21_X1 port map( B1 => n5462, B2 => n1659, A => n1661, ZN => n4028)
                           ;
   U888 : NAND2_X1 port map( A1 => n1659, A2 => n6706, ZN => n1661);
   U889 : OAI21_X1 port map( B1 => n5465, B2 => n5898, A => n1662, ZN => n4027)
                           ;
   U890 : NAND2_X1 port map( A1 => n1659, A2 => n6705, ZN => n1662);
   U891 : OAI21_X1 port map( B1 => n5468, B2 => n1659, A => n1663, ZN => n4026)
                           ;
   U892 : NAND2_X1 port map( A1 => n1659, A2 => n6704, ZN => n1663);
   U893 : OAI21_X1 port map( B1 => n5471, B2 => n1659, A => n1664, ZN => n4025)
                           ;
   U894 : NAND2_X1 port map( A1 => n5900, A2 => n6703, ZN => n1664);
   U895 : OAI21_X1 port map( B1 => n5474, B2 => n5898, A => n1665, ZN => n4024)
                           ;
   U896 : NAND2_X1 port map( A1 => n5900, A2 => n6702, ZN => n1665);
   U897 : OAI21_X1 port map( B1 => n5477, B2 => n5898, A => n1666, ZN => n4023)
                           ;
   U898 : NAND2_X1 port map( A1 => n1659, A2 => n6701, ZN => n1666);
   U899 : OAI21_X1 port map( B1 => n5480, B2 => n5898, A => n1667, ZN => n4022)
                           ;
   U900 : NAND2_X1 port map( A1 => n1659, A2 => n6700, ZN => n1667);
   U901 : OAI21_X1 port map( B1 => n6067, B2 => n5898, A => n1668, ZN => n4021)
                           ;
   U902 : NAND2_X1 port map( A1 => n1659, A2 => n6699, ZN => n1668);
   U903 : OAI21_X1 port map( B1 => n5486, B2 => n5898, A => n1669, ZN => n4020)
                           ;
   U904 : NAND2_X1 port map( A1 => n1659, A2 => n6698, ZN => n1669);
   U905 : OAI21_X1 port map( B1 => n5489, B2 => n5898, A => n1670, ZN => n4019)
                           ;
   U906 : NAND2_X1 port map( A1 => n1659, A2 => n6697, ZN => n1670);
   U907 : OAI21_X1 port map( B1 => n5492, B2 => n5898, A => n1671, ZN => n4018)
                           ;
   U908 : NAND2_X1 port map( A1 => n1659, A2 => n6696, ZN => n1671);
   U909 : OAI21_X1 port map( B1 => n5495, B2 => n5898, A => n1672, ZN => n4017)
                           ;
   U910 : NAND2_X1 port map( A1 => n1659, A2 => n6695, ZN => n1672);
   U911 : OAI21_X1 port map( B1 => n5498, B2 => n5898, A => n1673, ZN => n4016)
                           ;
   U912 : NAND2_X1 port map( A1 => n1659, A2 => n6694, ZN => n1673);
   U913 : OAI21_X1 port map( B1 => n6073, B2 => n5898, A => n1674, ZN => n4015)
                           ;
   U914 : NAND2_X1 port map( A1 => n1659, A2 => n6693, ZN => n1674);
   U915 : OAI21_X1 port map( B1 => n5504, B2 => n5900, A => n1675, ZN => n4014)
                           ;
   U916 : NAND2_X1 port map( A1 => n1659, A2 => n6692, ZN => n1675);
   U917 : OAI21_X1 port map( B1 => n6075, B2 => n5898, A => n1676, ZN => n4013)
                           ;
   U918 : NAND2_X1 port map( A1 => n5898, A2 => n6691, ZN => n1676);
   U919 : OAI21_X1 port map( B1 => n5509, B2 => n5900, A => n1677, ZN => n4012)
                           ;
   U920 : NAND2_X1 port map( A1 => n5900, A2 => n6690, ZN => n1677);
   U921 : OAI21_X1 port map( B1 => n5513, B2 => n5898, A => n1678, ZN => n4011)
                           ;
   U922 : NAND2_X1 port map( A1 => n5900, A2 => n6689, ZN => n1678);
   U923 : OAI21_X1 port map( B1 => n5516, B2 => n5900, A => n1679, ZN => n4010)
                           ;
   U924 : NAND2_X1 port map( A1 => n5900, A2 => n6688, ZN => n1679);
   U925 : OAI21_X1 port map( B1 => n5519, B2 => n5898, A => n1680, ZN => n4009)
                           ;
   U926 : NAND2_X1 port map( A1 => n5900, A2 => n6687, ZN => n1680);
   U927 : OAI21_X1 port map( B1 => n5522, B2 => n5900, A => n1681, ZN => n4008)
                           ;
   U928 : NAND2_X1 port map( A1 => n5900, A2 => n6686, ZN => n1681);
   U929 : OAI21_X1 port map( B1 => n6081, B2 => n5898, A => n1682, ZN => n4007)
                           ;
   U930 : NAND2_X1 port map( A1 => n5900, A2 => n6685, ZN => n1682);
   U931 : OAI21_X1 port map( B1 => n5528, B2 => n5900, A => n1683, ZN => n4006)
                           ;
   U932 : NAND2_X1 port map( A1 => n5900, A2 => n6684, ZN => n1683);
   U933 : OAI21_X1 port map( B1 => n5531, B2 => n5898, A => n1684, ZN => n4005)
                           ;
   U934 : NAND2_X1 port map( A1 => n1659, A2 => n6683, ZN => n1684);
   U935 : OAI21_X1 port map( B1 => n5534, B2 => n5900, A => n1685, ZN => n4004)
                           ;
   U936 : NAND2_X1 port map( A1 => n1659, A2 => n6682, ZN => n1685);
   U937 : OAI21_X1 port map( B1 => n5537, B2 => n5898, A => n1686, ZN => n4003)
                           ;
   U938 : NAND2_X1 port map( A1 => n1659, A2 => n6681, ZN => n1686);
   U939 : OAI21_X1 port map( B1 => n5540, B2 => n5900, A => n1687, ZN => n4002)
                           ;
   U940 : NAND2_X1 port map( A1 => n1659, A2 => n6680, ZN => n1687);
   U941 : OAI21_X1 port map( B1 => n5543, B2 => n5900, A => n1688, ZN => n4001)
                           ;
   U942 : NAND2_X1 port map( A1 => n5900, A2 => n6679, ZN => n1688);
   U943 : OAI21_X1 port map( B1 => n5546, B2 => n5900, A => n1689, ZN => n4000)
                           ;
   U944 : NAND2_X1 port map( A1 => n1659, A2 => n6678, ZN => n1689);
   U945 : OAI21_X1 port map( B1 => n5549, B2 => n5900, A => n1690, ZN => n3999)
                           ;
   U946 : NAND2_X1 port map( A1 => n1659, A2 => n6677, ZN => n1690);
   U947 : OAI21_X1 port map( B1 => n5552, B2 => n1659, A => n1691, ZN => n3998)
                           ;
   U948 : NAND2_X1 port map( A1 => n5898, A2 => n6676, ZN => n1691);
   U949 : NAND2_X1 port map( A1 => n1692, A2 => n1555, ZN => n1659);
   U950 : OAI21_X1 port map( B1 => n5459, B2 => n5890, A => n1694, ZN => n3918)
                           ;
   U951 : NAND2_X1 port map( A1 => n5894, A2 => n7115, ZN => n1694);
   U952 : OAI21_X1 port map( B1 => n5462, B2 => n1693, A => n1695, ZN => n3917)
                           ;
   U953 : NAND2_X1 port map( A1 => n5894, A2 => n7114, ZN => n1695);
   U954 : OAI21_X1 port map( B1 => n5465, B2 => n5894, A => n1696, ZN => n3916)
                           ;
   U955 : NAND2_X1 port map( A1 => n5894, A2 => n7113, ZN => n1696);
   U956 : OAI21_X1 port map( B1 => n5468, B2 => n1693, A => n1697, ZN => n3915)
                           ;
   U957 : NAND2_X1 port map( A1 => n5894, A2 => n7112, ZN => n1697);
   U958 : OAI21_X1 port map( B1 => n5471, B2 => n1693, A => n1698, ZN => n3914)
                           ;
   U959 : NAND2_X1 port map( A1 => n5890, A2 => n7111, ZN => n1698);
   U960 : OAI21_X1 port map( B1 => n5474, B2 => n5894, A => n1699, ZN => n3913)
                           ;
   U961 : NAND2_X1 port map( A1 => n5890, A2 => n7110, ZN => n1699);
   U962 : OAI21_X1 port map( B1 => n5477, B2 => n5890, A => n1700, ZN => n3912)
                           ;
   U963 : NAND2_X1 port map( A1 => n5890, A2 => n7109, ZN => n1700);
   U964 : OAI21_X1 port map( B1 => n5480, B2 => n5890, A => n1701, ZN => n3911)
                           ;
   U965 : NAND2_X1 port map( A1 => n1693, A2 => n7108, ZN => n1701);
   U966 : OAI21_X1 port map( B1 => n6067, B2 => n5894, A => n1702, ZN => n3910)
                           ;
   U967 : NAND2_X1 port map( A1 => n1693, A2 => n7107, ZN => n1702);
   U968 : OAI21_X1 port map( B1 => n5486, B2 => n5890, A => n1703, ZN => n3909)
                           ;
   U969 : NAND2_X1 port map( A1 => n1693, A2 => n7106, ZN => n1703);
   U970 : OAI21_X1 port map( B1 => n5489, B2 => n5894, A => n1704, ZN => n3908)
                           ;
   U971 : NAND2_X1 port map( A1 => n1693, A2 => n7105, ZN => n1704);
   U972 : OAI21_X1 port map( B1 => n5492, B2 => n5890, A => n1705, ZN => n3907)
                           ;
   U973 : NAND2_X1 port map( A1 => n5890, A2 => n7104, ZN => n1705);
   U974 : OAI21_X1 port map( B1 => n5495, B2 => n5894, A => n1706, ZN => n3906)
                           ;
   U975 : NAND2_X1 port map( A1 => n5894, A2 => n7103, ZN => n1706);
   U976 : OAI21_X1 port map( B1 => n5498, B2 => n5894, A => n1707, ZN => n3905)
                           ;
   U977 : NAND2_X1 port map( A1 => n5890, A2 => n7102, ZN => n1707);
   U978 : OAI21_X1 port map( B1 => n6073, B2 => n5890, A => n1708, ZN => n3904)
                           ;
   U979 : NAND2_X1 port map( A1 => n1693, A2 => n7101, ZN => n1708);
   U980 : OAI21_X1 port map( B1 => n5504, B2 => n1693, A => n1709, ZN => n3903)
                           ;
   U981 : NAND2_X1 port map( A1 => n1693, A2 => n7100, ZN => n1709);
   U982 : OAI21_X1 port map( B1 => n6075, B2 => n1693, A => n1710, ZN => n3902)
                           ;
   U983 : NAND2_X1 port map( A1 => n5890, A2 => n7099, ZN => n1710);
   U984 : OAI21_X1 port map( B1 => n5509, B2 => n1693, A => n1711, ZN => n3901)
                           ;
   U985 : NAND2_X1 port map( A1 => n5890, A2 => n7098, ZN => n1711);
   U986 : OAI21_X1 port map( B1 => n5513, B2 => n1693, A => n1712, ZN => n3900)
                           ;
   U987 : NAND2_X1 port map( A1 => n5890, A2 => n7097, ZN => n1712);
   U988 : OAI21_X1 port map( B1 => n5516, B2 => n1693, A => n1713, ZN => n3899)
                           ;
   U989 : NAND2_X1 port map( A1 => n5890, A2 => n7096, ZN => n1713);
   U990 : OAI21_X1 port map( B1 => n5519, B2 => n1693, A => n1714, ZN => n3898)
                           ;
   U991 : NAND2_X1 port map( A1 => n5890, A2 => n7095, ZN => n1714);
   U992 : OAI21_X1 port map( B1 => n5522, B2 => n1693, A => n1715, ZN => n3897)
                           ;
   U993 : NAND2_X1 port map( A1 => n5890, A2 => n7094, ZN => n1715);
   U994 : OAI21_X1 port map( B1 => n6081, B2 => n1693, A => n1716, ZN => n3896)
                           ;
   U995 : NAND2_X1 port map( A1 => n5890, A2 => n7093, ZN => n1716);
   U996 : OAI21_X1 port map( B1 => n5528, B2 => n1693, A => n1717, ZN => n3895)
                           ;
   U997 : NAND2_X1 port map( A1 => n5890, A2 => n7092, ZN => n1717);
   U998 : OAI21_X1 port map( B1 => n5531, B2 => n1693, A => n1718, ZN => n3894)
                           ;
   U999 : NAND2_X1 port map( A1 => n5894, A2 => n7091, ZN => n1718);
   U1000 : OAI21_X1 port map( B1 => n5534, B2 => n1693, A => n1719, ZN => n3893
                           );
   U1001 : NAND2_X1 port map( A1 => n5894, A2 => n7090, ZN => n1719);
   U1002 : OAI21_X1 port map( B1 => n5537, B2 => n1693, A => n1720, ZN => n3892
                           );
   U1003 : NAND2_X1 port map( A1 => n5894, A2 => n7089, ZN => n1720);
   U1004 : OAI21_X1 port map( B1 => n5540, B2 => n5894, A => n1721, ZN => n3891
                           );
   U1005 : NAND2_X1 port map( A1 => n5894, A2 => n7088, ZN => n1721);
   U1006 : OAI21_X1 port map( B1 => n5543, B2 => n5894, A => n1722, ZN => n3890
                           );
   U1007 : NAND2_X1 port map( A1 => n5890, A2 => n7087, ZN => n1722);
   U1008 : OAI21_X1 port map( B1 => n5546, B2 => n5894, A => n1723, ZN => n3889
                           );
   U1009 : NAND2_X1 port map( A1 => n1693, A2 => n7086, ZN => n1723);
   U1010 : OAI21_X1 port map( B1 => n5549, B2 => n5894, A => n1724, ZN => n3888
                           );
   U1011 : NAND2_X1 port map( A1 => n1693, A2 => n7085, ZN => n1724);
   U1012 : OAI21_X1 port map( B1 => n5552, B2 => n1693, A => n1725, ZN => n3887
                           );
   U1013 : NAND2_X1 port map( A1 => n5894, A2 => n7084, ZN => n1725);
   U1014 : NAND2_X1 port map( A1 => n1692, A2 => n1658, ZN => n1693);
   U1015 : OAI21_X1 port map( B1 => n5459, B2 => n5886, A => n1727, ZN => n3886
                           );
   U1016 : NAND2_X1 port map( A1 => n1726, A2 => n6859, ZN => n1727);
   U1017 : OAI21_X1 port map( B1 => n5462, B2 => n5887, A => n1728, ZN => n3885
                           );
   U1018 : NAND2_X1 port map( A1 => n1726, A2 => n6858, ZN => n1728);
   U1019 : OAI21_X1 port map( B1 => n5465, B2 => n5886, A => n1729, ZN => n3884
                           );
   U1020 : NAND2_X1 port map( A1 => n1726, A2 => n6857, ZN => n1729);
   U1021 : OAI21_X1 port map( B1 => n5468, B2 => n5886, A => n1730, ZN => n3883
                           );
   U1022 : NAND2_X1 port map( A1 => n1726, A2 => n6856, ZN => n1730);
   U1023 : OAI21_X1 port map( B1 => n5471, B2 => n5887, A => n1731, ZN => n3882
                           );
   U1024 : NAND2_X1 port map( A1 => n1726, A2 => n6855, ZN => n1731);
   U1025 : OAI21_X1 port map( B1 => n5474, B2 => n5886, A => n1732, ZN => n3881
                           );
   U1026 : NAND2_X1 port map( A1 => n1726, A2 => n6854, ZN => n1732);
   U1027 : OAI21_X1 port map( B1 => n5477, B2 => n5886, A => n1733, ZN => n3880
                           );
   U1028 : NAND2_X1 port map( A1 => n1726, A2 => n6853, ZN => n1733);
   U1029 : OAI21_X1 port map( B1 => n5480, B2 => n5886, A => n1734, ZN => n3879
                           );
   U1030 : NAND2_X1 port map( A1 => n5887, A2 => n6852, ZN => n1734);
   U1031 : OAI21_X1 port map( B1 => n6067, B2 => n5886, A => n1735, ZN => n3878
                           );
   U1032 : NAND2_X1 port map( A1 => n5886, A2 => n6851, ZN => n1735);
   U1033 : OAI21_X1 port map( B1 => n5486, B2 => n5886, A => n1736, ZN => n3877
                           );
   U1034 : NAND2_X1 port map( A1 => n5887, A2 => n6850, ZN => n1736);
   U1035 : OAI21_X1 port map( B1 => n5489, B2 => n5886, A => n1737, ZN => n3876
                           );
   U1036 : NAND2_X1 port map( A1 => n5886, A2 => n6849, ZN => n1737);
   U1037 : OAI21_X1 port map( B1 => n5492, B2 => n5886, A => n1738, ZN => n3875
                           );
   U1038 : NAND2_X1 port map( A1 => n5887, A2 => n6848, ZN => n1738);
   U1039 : OAI21_X1 port map( B1 => n5495, B2 => n5886, A => n1739, ZN => n3874
                           );
   U1040 : NAND2_X1 port map( A1 => n5886, A2 => n6847, ZN => n1739);
   U1041 : OAI21_X1 port map( B1 => n5498, B2 => n5886, A => n1740, ZN => n3873
                           );
   U1042 : NAND2_X1 port map( A1 => n1726, A2 => n6846, ZN => n1740);
   U1043 : OAI21_X1 port map( B1 => n6073, B2 => n5886, A => n1741, ZN => n3872
                           );
   U1044 : NAND2_X1 port map( A1 => n5887, A2 => n6845, ZN => n1741);
   U1045 : OAI21_X1 port map( B1 => n5504, B2 => n5887, A => n1742, ZN => n3871
                           );
   U1046 : NAND2_X1 port map( A1 => n5886, A2 => n6844, ZN => n1742);
   U1047 : OAI21_X1 port map( B1 => n6075, B2 => n5887, A => n1743, ZN => n3870
                           );
   U1048 : NAND2_X1 port map( A1 => n1726, A2 => n6843, ZN => n1743);
   U1049 : OAI21_X1 port map( B1 => n5459, B2 => n5880, A => n1745, ZN => n3869
                           );
   U1050 : NAND2_X1 port map( A1 => n2830, A2 => n1744, ZN => n1745);
   U1051 : OAI21_X1 port map( B1 => n5462, B2 => n1744, A => n1746, ZN => n3868
                           );
   U1052 : NAND2_X1 port map( A1 => n2829, A2 => n5882, ZN => n1746);
   U1053 : OAI21_X1 port map( B1 => n5465, B2 => n5880, A => n1747, ZN => n3867
                           );
   U1054 : NAND2_X1 port map( A1 => n2828, A2 => n1744, ZN => n1747);
   U1055 : OAI21_X1 port map( B1 => n5468, B2 => n1744, A => n1748, ZN => n3866
                           );
   U1056 : NAND2_X1 port map( A1 => n2827, A2 => n5880, ZN => n1748);
   U1057 : OAI21_X1 port map( B1 => n5471, B2 => n1744, A => n1749, ZN => n3865
                           );
   U1058 : NAND2_X1 port map( A1 => n2826, A2 => n5882, ZN => n1749);
   U1059 : OAI21_X1 port map( B1 => n5474, B2 => n5880, A => n1750, ZN => n3864
                           );
   U1060 : NAND2_X1 port map( A1 => n2825, A2 => n1744, ZN => n1750);
   U1061 : OAI21_X1 port map( B1 => n5477, B2 => n5880, A => n1751, ZN => n3863
                           );
   U1062 : NAND2_X1 port map( A1 => n2824, A2 => n1744, ZN => n1751);
   U1063 : OAI21_X1 port map( B1 => n5480, B2 => n5880, A => n1752, ZN => n3862
                           );
   U1064 : NAND2_X1 port map( A1 => n2823, A2 => n5882, ZN => n1752);
   U1065 : OAI21_X1 port map( B1 => n6067, B2 => n5880, A => n1753, ZN => n3861
                           );
   U1066 : NAND2_X1 port map( A1 => n2822, A2 => n1744, ZN => n1753);
   U1067 : OAI21_X1 port map( B1 => n5486, B2 => n5880, A => n1754, ZN => n3860
                           );
   U1068 : NAND2_X1 port map( A1 => n2821, A2 => n1744, ZN => n1754);
   U1069 : OAI21_X1 port map( B1 => n5489, B2 => n5880, A => n1755, ZN => n3859
                           );
   U1070 : NAND2_X1 port map( A1 => n2820, A2 => n5880, ZN => n1755);
   U1071 : OAI21_X1 port map( B1 => n5492, B2 => n5880, A => n1756, ZN => n3858
                           );
   U1072 : NAND2_X1 port map( A1 => n2819, A2 => n5882, ZN => n1756);
   U1073 : OAI21_X1 port map( B1 => n5495, B2 => n5880, A => n1757, ZN => n3857
                           );
   U1074 : NAND2_X1 port map( A1 => n2818, A2 => n5882, ZN => n1757);
   U1075 : OAI21_X1 port map( B1 => n5498, B2 => n5880, A => n1758, ZN => n3856
                           );
   U1076 : NAND2_X1 port map( A1 => n2817, A2 => n5882, ZN => n1758);
   U1077 : OAI21_X1 port map( B1 => n6073, B2 => n5880, A => n1759, ZN => n3855
                           );
   U1078 : NAND2_X1 port map( A1 => n2816, A2 => n1744, ZN => n1759);
   U1079 : OAI21_X1 port map( B1 => n5504, B2 => n5882, A => n1760, ZN => n3854
                           );
   U1080 : NAND2_X1 port map( A1 => n2815, A2 => n5882, ZN => n1760);
   U1081 : OAI21_X1 port map( B1 => n6075, B2 => n5880, A => n1761, ZN => n3853
                           );
   U1082 : NAND2_X1 port map( A1 => n2814, A2 => n1744, ZN => n1761);
   U1083 : OAI21_X1 port map( B1 => n5509, B2 => n5882, A => n1762, ZN => n3852
                           );
   U1084 : NAND2_X1 port map( A1 => n2813, A2 => n5882, ZN => n1762);
   U1085 : OAI21_X1 port map( B1 => n5513, B2 => n5880, A => n1763, ZN => n3851
                           );
   U1086 : NAND2_X1 port map( A1 => n2812, A2 => n1744, ZN => n1763);
   U1087 : OAI21_X1 port map( B1 => n5516, B2 => n5882, A => n1764, ZN => n3850
                           );
   U1088 : NAND2_X1 port map( A1 => n2811, A2 => n1744, ZN => n1764);
   U1089 : OAI21_X1 port map( B1 => n5519, B2 => n5880, A => n1765, ZN => n3849
                           );
   U1090 : NAND2_X1 port map( A1 => n2810, A2 => n5882, ZN => n1765);
   U1091 : OAI21_X1 port map( B1 => n5522, B2 => n5882, A => n1766, ZN => n3848
                           );
   U1092 : NAND2_X1 port map( A1 => n2809, A2 => n5882, ZN => n1766);
   U1093 : OAI21_X1 port map( B1 => n6081, B2 => n5880, A => n1767, ZN => n3847
                           );
   U1094 : NAND2_X1 port map( A1 => n2808, A2 => n5882, ZN => n1767);
   U1095 : OAI21_X1 port map( B1 => n5528, B2 => n5882, A => n1768, ZN => n3846
                           );
   U1096 : NAND2_X1 port map( A1 => n2807, A2 => n5880, ZN => n1768);
   U1097 : OAI21_X1 port map( B1 => n5531, B2 => n5880, A => n1769, ZN => n3845
                           );
   U1098 : NAND2_X1 port map( A1 => n1744, A2 => n6675, ZN => n1769);
   U1099 : OAI21_X1 port map( B1 => n5534, B2 => n1744, A => n1770, ZN => n3844
                           );
   U1100 : NAND2_X1 port map( A1 => n1744, A2 => n6674, ZN => n1770);
   U1101 : OAI21_X1 port map( B1 => n5537, B2 => n1744, A => n1771, ZN => n3843
                           );
   U1102 : NAND2_X1 port map( A1 => n1744, A2 => n6673, ZN => n1771);
   U1103 : OAI21_X1 port map( B1 => n5540, B2 => n5882, A => n1772, ZN => n3842
                           );
   U1104 : NAND2_X1 port map( A1 => n1744, A2 => n6672, ZN => n1772);
   U1105 : OAI21_X1 port map( B1 => n5543, B2 => n5882, A => n1773, ZN => n3841
                           );
   U1106 : NAND2_X1 port map( A1 => n1744, A2 => n6671, ZN => n1773);
   U1107 : OAI21_X1 port map( B1 => n5546, B2 => n5882, A => n1774, ZN => n3840
                           );
   U1108 : NAND2_X1 port map( A1 => n1744, A2 => n6670, ZN => n1774);
   U1109 : OAI21_X1 port map( B1 => n5549, B2 => n5882, A => n1775, ZN => n3839
                           );
   U1110 : NAND2_X1 port map( A1 => n1744, A2 => n6669, ZN => n1775);
   U1111 : OAI21_X1 port map( B1 => n5552, B2 => n1744, A => n1776, ZN => n3838
                           );
   U1112 : NAND2_X1 port map( A1 => n1744, A2 => n6668, ZN => n1776);
   U1113 : NAND2_X1 port map( A1 => n1777, A2 => n1778, ZN => n1744);
   U1114 : OAI21_X1 port map( B1 => n5459, B2 => n1779, A => n1780, ZN => n3837
                           );
   U1115 : NAND2_X1 port map( A1 => n5871, A2 => n6742, ZN => n1780);
   U1116 : OAI21_X1 port map( B1 => n5462, B2 => n5873, A => n1781, ZN => n3836
                           );
   U1117 : NAND2_X1 port map( A1 => n5871, A2 => n6741, ZN => n1781);
   U1118 : OAI21_X1 port map( B1 => n5465, B2 => n1779, A => n1782, ZN => n3835
                           );
   U1119 : NAND2_X1 port map( A1 => n5871, A2 => n6740, ZN => n1782);
   U1120 : OAI21_X1 port map( B1 => n5468, B2 => n5873, A => n1783, ZN => n3834
                           );
   U1121 : NAND2_X1 port map( A1 => n5871, A2 => n6739, ZN => n1783);
   U1122 : OAI21_X1 port map( B1 => n5471, B2 => n5873, A => n1784, ZN => n3833
                           );
   U1123 : NAND2_X1 port map( A1 => n5871, A2 => n6738, ZN => n1784);
   U1124 : OAI21_X1 port map( B1 => n5474, B2 => n1779, A => n1785, ZN => n3832
                           );
   U1125 : NAND2_X1 port map( A1 => n5873, A2 => n6737, ZN => n1785);
   U1126 : OAI21_X1 port map( B1 => n5477, B2 => n1779, A => n1786, ZN => n3831
                           );
   U1127 : NAND2_X1 port map( A1 => n5871, A2 => n6736, ZN => n1786);
   U1128 : OAI21_X1 port map( B1 => n5480, B2 => n1779, A => n1787, ZN => n3830
                           );
   U1129 : NAND2_X1 port map( A1 => n5873, A2 => n6735, ZN => n1787);
   U1130 : OAI21_X1 port map( B1 => n6067, B2 => n1779, A => n1788, ZN => n3829
                           );
   U1131 : NAND2_X1 port map( A1 => n5873, A2 => n6734, ZN => n1788);
   U1132 : OAI21_X1 port map( B1 => n5486, B2 => n1779, A => n1789, ZN => n3828
                           );
   U1133 : NAND2_X1 port map( A1 => n5873, A2 => n6733, ZN => n1789);
   U1134 : OAI21_X1 port map( B1 => n5489, B2 => n1779, A => n1790, ZN => n3827
                           );
   U1135 : NAND2_X1 port map( A1 => n5873, A2 => n6732, ZN => n1790);
   U1136 : OAI21_X1 port map( B1 => n5492, B2 => n1779, A => n1791, ZN => n3826
                           );
   U1137 : NAND2_X1 port map( A1 => n5873, A2 => n6731, ZN => n1791);
   U1138 : OAI21_X1 port map( B1 => n5495, B2 => n1779, A => n1792, ZN => n3825
                           );
   U1139 : NAND2_X1 port map( A1 => n5873, A2 => n6730, ZN => n1792);
   U1140 : OAI21_X1 port map( B1 => n5498, B2 => n1779, A => n1793, ZN => n3824
                           );
   U1141 : NAND2_X1 port map( A1 => n5873, A2 => n6729, ZN => n1793);
   U1142 : OAI21_X1 port map( B1 => n6073, B2 => n1779, A => n1794, ZN => n3823
                           );
   U1143 : NAND2_X1 port map( A1 => n5873, A2 => n6728, ZN => n1794);
   U1144 : OAI21_X1 port map( B1 => n5504, B2 => n1779, A => n1795, ZN => n3822
                           );
   U1145 : NAND2_X1 port map( A1 => n5873, A2 => n6727, ZN => n1795);
   U1146 : OAI21_X1 port map( B1 => n5506, B2 => n1779, A => n1796, ZN => n3821
                           );
   U1147 : NAND2_X1 port map( A1 => n5871, A2 => n6726, ZN => n1796);
   U1148 : OAI21_X1 port map( B1 => n5509, B2 => n5873, A => n1797, ZN => n3820
                           );
   U1149 : NAND2_X1 port map( A1 => n5873, A2 => n6725, ZN => n1797);
   U1150 : OAI21_X1 port map( B1 => n5513, B2 => n1779, A => n1798, ZN => n3819
                           );
   U1151 : NAND2_X1 port map( A1 => n5873, A2 => n6724, ZN => n1798);
   U1152 : OAI21_X1 port map( B1 => n5516, B2 => n5873, A => n1799, ZN => n3818
                           );
   U1153 : NAND2_X1 port map( A1 => n5871, A2 => n6723, ZN => n1799);
   U1154 : OAI21_X1 port map( B1 => n5519, B2 => n1779, A => n1800, ZN => n3817
                           );
   U1155 : NAND2_X1 port map( A1 => n5873, A2 => n6722, ZN => n1800);
   U1156 : OAI21_X1 port map( B1 => n5522, B2 => n5871, A => n1801, ZN => n3816
                           );
   U1157 : NAND2_X1 port map( A1 => n5871, A2 => n6721, ZN => n1801);
   U1158 : OAI21_X1 port map( B1 => n6081, B2 => n5873, A => n1802, ZN => n3815
                           );
   U1159 : NAND2_X1 port map( A1 => n5871, A2 => n6720, ZN => n1802);
   U1160 : OAI21_X1 port map( B1 => n5528, B2 => n1779, A => n1803, ZN => n3814
                           );
   U1161 : NAND2_X1 port map( A1 => n5871, A2 => n6719, ZN => n1803);
   U1162 : OAI21_X1 port map( B1 => n5531, B2 => n1779, A => n1804, ZN => n3813
                           );
   U1163 : NAND2_X1 port map( A1 => n5871, A2 => n6718, ZN => n1804);
   U1164 : OAI21_X1 port map( B1 => n5534, B2 => n1779, A => n1805, ZN => n3812
                           );
   U1165 : NAND2_X1 port map( A1 => n5871, A2 => n6717, ZN => n1805);
   U1166 : OAI21_X1 port map( B1 => n5537, B2 => n1779, A => n1806, ZN => n3811
                           );
   U1167 : NAND2_X1 port map( A1 => n5871, A2 => n6716, ZN => n1806);
   U1168 : OAI21_X1 port map( B1 => n5540, B2 => n1779, A => n1807, ZN => n3810
                           );
   U1169 : NAND2_X1 port map( A1 => n5871, A2 => n6715, ZN => n1807);
   U1170 : OAI21_X1 port map( B1 => n5543, B2 => n1779, A => n1808, ZN => n3809
                           );
   U1171 : NAND2_X1 port map( A1 => n5871, A2 => n6714, ZN => n1808);
   U1172 : OAI21_X1 port map( B1 => n5546, B2 => n1779, A => n1809, ZN => n3808
                           );
   U1173 : NAND2_X1 port map( A1 => n5871, A2 => n6713, ZN => n1809);
   U1174 : OAI21_X1 port map( B1 => n5549, B2 => n1779, A => n1810, ZN => n3807
                           );
   U1175 : NAND2_X1 port map( A1 => n5871, A2 => n6712, ZN => n1810);
   U1176 : OAI21_X1 port map( B1 => n5552, B2 => n5873, A => n1811, ZN => n3806
                           );
   U1177 : NAND2_X1 port map( A1 => n5871, A2 => n6711, ZN => n1811);
   U1178 : NAND2_X1 port map( A1 => n1812, A2 => n1777, ZN => n1779);
   U1179 : OAI21_X1 port map( B1 => n5509, B2 => n5887, A => n1813, ZN => n3805
                           );
   U1180 : NAND2_X1 port map( A1 => n1726, A2 => n6842, ZN => n1813);
   U1181 : OAI21_X1 port map( B1 => n5513, B2 => n5887, A => n1814, ZN => n3804
                           );
   U1182 : NAND2_X1 port map( A1 => n1726, A2 => n6841, ZN => n1814);
   U1183 : OAI21_X1 port map( B1 => n5516, B2 => n5887, A => n1815, ZN => n3803
                           );
   U1184 : NAND2_X1 port map( A1 => n1726, A2 => n6840, ZN => n1815);
   U1185 : OAI21_X1 port map( B1 => n5519, B2 => n5887, A => n1816, ZN => n3802
                           );
   U1186 : NAND2_X1 port map( A1 => n1726, A2 => n6839, ZN => n1816);
   U1187 : OAI21_X1 port map( B1 => n5522, B2 => n5887, A => n1817, ZN => n3801
                           );
   U1188 : NAND2_X1 port map( A1 => n1726, A2 => n6838, ZN => n1817);
   U1189 : OAI21_X1 port map( B1 => n6081, B2 => n5887, A => n1818, ZN => n3800
                           );
   U1190 : NAND2_X1 port map( A1 => n1726, A2 => n6837, ZN => n1818);
   U1191 : OAI21_X1 port map( B1 => n5528, B2 => n5887, A => n1819, ZN => n3799
                           );
   U1192 : NAND2_X1 port map( A1 => n1726, A2 => n6836, ZN => n1819);
   U1193 : OAI21_X1 port map( B1 => n5531, B2 => n5887, A => n1820, ZN => n3798
                           );
   U1194 : NAND2_X1 port map( A1 => n1726, A2 => n6835, ZN => n1820);
   U1195 : OAI21_X1 port map( B1 => n5534, B2 => n5887, A => n1821, ZN => n3797
                           );
   U1196 : NAND2_X1 port map( A1 => n1726, A2 => n6834, ZN => n1821);
   U1197 : OAI21_X1 port map( B1 => n5537, B2 => n5887, A => n1822, ZN => n3796
                           );
   U1198 : NAND2_X1 port map( A1 => n1726, A2 => n6833, ZN => n1822);
   U1199 : OAI21_X1 port map( B1 => n5540, B2 => n5887, A => n1823, ZN => n3795
                           );
   U1200 : NAND2_X1 port map( A1 => n1726, A2 => n6832, ZN => n1823);
   U1201 : OAI21_X1 port map( B1 => n5543, B2 => n5886, A => n1824, ZN => n3794
                           );
   U1202 : NAND2_X1 port map( A1 => n1726, A2 => n6831, ZN => n1824);
   U1203 : OAI21_X1 port map( B1 => n5546, B2 => n5887, A => n1825, ZN => n3793
                           );
   U1204 : NAND2_X1 port map( A1 => n1726, A2 => n6830, ZN => n1825);
   U1205 : OAI21_X1 port map( B1 => n5549, B2 => n5886, A => n1826, ZN => n3792
                           );
   U1206 : NAND2_X1 port map( A1 => n1726, A2 => n6829, ZN => n1826);
   U1207 : OAI21_X1 port map( B1 => n5552, B2 => n5886, A => n1827, ZN => n3791
                           );
   U1208 : NAND2_X1 port map( A1 => n1726, A2 => n6828, ZN => n1827);
   U1209 : NAND2_X1 port map( A1 => n1692, A2 => n1624, ZN => n1726);
   U1210 : OAI21_X1 port map( B1 => n5459, B2 => n5868, A => n1829, ZN => n3790
                           );
   U1211 : NAND2_X1 port map( A1 => n1828, A2 => n6987, ZN => n1829);
   U1212 : OAI21_X1 port map( B1 => n5462, B2 => n5869, A => n1830, ZN => n3789
                           );
   U1213 : NAND2_X1 port map( A1 => n1828, A2 => n6986, ZN => n1830);
   U1214 : OAI21_X1 port map( B1 => n5465, B2 => n5868, A => n1831, ZN => n3788
                           );
   U1215 : NAND2_X1 port map( A1 => n1828, A2 => n6985, ZN => n1831);
   U1216 : OAI21_X1 port map( B1 => n5468, B2 => n5868, A => n1832, ZN => n3787
                           );
   U1217 : NAND2_X1 port map( A1 => n1828, A2 => n6984, ZN => n1832);
   U1218 : OAI21_X1 port map( B1 => n5471, B2 => n5869, A => n1833, ZN => n3786
                           );
   U1219 : NAND2_X1 port map( A1 => n1828, A2 => n6983, ZN => n1833);
   U1220 : OAI21_X1 port map( B1 => n5474, B2 => n5868, A => n1834, ZN => n3785
                           );
   U1221 : NAND2_X1 port map( A1 => n1828, A2 => n6982, ZN => n1834);
   U1222 : OAI21_X1 port map( B1 => n5477, B2 => n5868, A => n1835, ZN => n3784
                           );
   U1223 : NAND2_X1 port map( A1 => n1828, A2 => n6981, ZN => n1835);
   U1224 : OAI21_X1 port map( B1 => n5480, B2 => n5868, A => n1836, ZN => n3783
                           );
   U1225 : NAND2_X1 port map( A1 => n5869, A2 => n6980, ZN => n1836);
   U1226 : OAI21_X1 port map( B1 => n6067, B2 => n5868, A => n1837, ZN => n3782
                           );
   U1227 : NAND2_X1 port map( A1 => n5868, A2 => n6979, ZN => n1837);
   U1228 : OAI21_X1 port map( B1 => n5486, B2 => n5868, A => n1838, ZN => n3781
                           );
   U1229 : NAND2_X1 port map( A1 => n5869, A2 => n6978, ZN => n1838);
   U1230 : OAI21_X1 port map( B1 => n5489, B2 => n5868, A => n1839, ZN => n3780
                           );
   U1231 : NAND2_X1 port map( A1 => n5868, A2 => n6977, ZN => n1839);
   U1232 : OAI21_X1 port map( B1 => n5492, B2 => n5868, A => n1840, ZN => n3779
                           );
   U1233 : NAND2_X1 port map( A1 => n5869, A2 => n6976, ZN => n1840);
   U1234 : OAI21_X1 port map( B1 => n5495, B2 => n5868, A => n1841, ZN => n3778
                           );
   U1235 : NAND2_X1 port map( A1 => n5868, A2 => n6975, ZN => n1841);
   U1236 : OAI21_X1 port map( B1 => n5498, B2 => n5868, A => n1842, ZN => n3777
                           );
   U1237 : NAND2_X1 port map( A1 => n1828, A2 => n6974, ZN => n1842);
   U1238 : OAI21_X1 port map( B1 => n6073, B2 => n5868, A => n1843, ZN => n3776
                           );
   U1239 : NAND2_X1 port map( A1 => n5869, A2 => n6973, ZN => n1843);
   U1240 : OAI21_X1 port map( B1 => n5504, B2 => n5869, A => n1844, ZN => n3775
                           );
   U1241 : NAND2_X1 port map( A1 => n5868, A2 => n6972, ZN => n1844);
   U1242 : OAI21_X1 port map( B1 => n5506, B2 => n5869, A => n1845, ZN => n3774
                           );
   U1243 : NAND2_X1 port map( A1 => n1828, A2 => n6971, ZN => n1845);
   U1244 : OAI21_X1 port map( B1 => n5552, B2 => n5864, A => n1847, ZN => n3773
                           );
   U1245 : NAND2_X1 port map( A1 => n321, A2 => n1846, ZN => n1847);
   U1246 : OAI21_X1 port map( B1 => n5549, B2 => n1846, A => n1848, ZN => n3772
                           );
   U1247 : NAND2_X1 port map( A1 => n322, A2 => n1846, ZN => n1848);
   U1248 : OAI21_X1 port map( B1 => n5546, B2 => n5863, A => n1849, ZN => n3771
                           );
   U1249 : NAND2_X1 port map( A1 => n323, A2 => n1846, ZN => n1849);
   U1250 : OAI21_X1 port map( B1 => n5543, B2 => n1846, A => n1850, ZN => n3770
                           );
   U1251 : NAND2_X1 port map( A1 => n324, A2 => n1846, ZN => n1850);
   U1252 : OAI21_X1 port map( B1 => n5540, B2 => n1846, A => n1851, ZN => n3769
                           );
   U1253 : NAND2_X1 port map( A1 => n325, A2 => n5864, ZN => n1851);
   U1254 : OAI21_X1 port map( B1 => n5537, B2 => n5864, A => n1852, ZN => n3768
                           );
   U1255 : NAND2_X1 port map( A1 => n326, A2 => n5864, ZN => n1852);
   U1256 : OAI21_X1 port map( B1 => n5534, B2 => n5863, A => n1853, ZN => n3767
                           );
   U1257 : NAND2_X1 port map( A1 => n327, A2 => n1846, ZN => n1853);
   U1258 : OAI21_X1 port map( B1 => n5531, B2 => n5864, A => n1854, ZN => n3766
                           );
   U1259 : NAND2_X1 port map( A1 => n328, A2 => n1846, ZN => n1854);
   U1260 : OAI21_X1 port map( B1 => n5528, B2 => n5863, A => n1855, ZN => n3765
                           );
   U1261 : NAND2_X1 port map( A1 => n329, A2 => n1846, ZN => n1855);
   U1262 : OAI21_X1 port map( B1 => n6081, B2 => n5864, A => n1856, ZN => n3764
                           );
   U1263 : NAND2_X1 port map( A1 => n330, A2 => n1846, ZN => n1856);
   U1264 : OAI21_X1 port map( B1 => n5522, B2 => n5863, A => n1857, ZN => n3763
                           );
   U1265 : NAND2_X1 port map( A1 => n331, A2 => n1846, ZN => n1857);
   U1266 : OAI21_X1 port map( B1 => n5519, B2 => n5864, A => n1858, ZN => n3762
                           );
   U1267 : NAND2_X1 port map( A1 => n332, A2 => n1846, ZN => n1858);
   U1268 : OAI21_X1 port map( B1 => n5516, B2 => n5863, A => n1859, ZN => n3761
                           );
   U1269 : NAND2_X1 port map( A1 => n333, A2 => n1846, ZN => n1859);
   U1270 : OAI21_X1 port map( B1 => n5513, B2 => n1846, A => n1860, ZN => n3760
                           );
   U1271 : NAND2_X1 port map( A1 => n334, A2 => n5864, ZN => n1860);
   U1272 : OAI21_X1 port map( B1 => n5509, B2 => n1846, A => n1861, ZN => n3759
                           );
   U1273 : NAND2_X1 port map( A1 => n335, A2 => n1846, ZN => n1861);
   U1274 : OAI21_X1 port map( B1 => n5506, B2 => n5863, A => n1862, ZN => n3758
                           );
   U1275 : NAND2_X1 port map( A1 => n336, A2 => n1846, ZN => n1862);
   U1276 : OAI21_X1 port map( B1 => n5504, B2 => n5863, A => n1863, ZN => n3757
                           );
   U1277 : NAND2_X1 port map( A1 => n337, A2 => n5863, ZN => n1863);
   U1278 : OAI21_X1 port map( B1 => n6073, B2 => n5863, A => n1864, ZN => n3756
                           );
   U1279 : NAND2_X1 port map( A1 => n338, A2 => n5864, ZN => n1864);
   U1280 : OAI21_X1 port map( B1 => n5498, B2 => n5863, A => n1865, ZN => n3755
                           );
   U1281 : NAND2_X1 port map( A1 => n339, A2 => n5864, ZN => n1865);
   U1282 : OAI21_X1 port map( B1 => n5495, B2 => n5863, A => n1866, ZN => n3754
                           );
   U1283 : NAND2_X1 port map( A1 => n340, A2 => n5864, ZN => n1866);
   U1284 : OAI21_X1 port map( B1 => n5492, B2 => n5863, A => n1867, ZN => n3753
                           );
   U1285 : NAND2_X1 port map( A1 => n341, A2 => n5864, ZN => n1867);
   U1286 : OAI21_X1 port map( B1 => n5489, B2 => n5863, A => n1868, ZN => n3752
                           );
   U1287 : NAND2_X1 port map( A1 => n342, A2 => n5864, ZN => n1868);
   U1288 : OAI21_X1 port map( B1 => n5486, B2 => n5863, A => n1869, ZN => n3751
                           );
   U1289 : NAND2_X1 port map( A1 => n343, A2 => n5864, ZN => n1869);
   U1290 : OAI21_X1 port map( B1 => n6067, B2 => n5863, A => n1870, ZN => n3750
                           );
   U1291 : NAND2_X1 port map( A1 => n344, A2 => n5864, ZN => n1870);
   U1292 : OAI21_X1 port map( B1 => n5480, B2 => n5863, A => n1871, ZN => n3749
                           );
   U1293 : NAND2_X1 port map( A1 => n345, A2 => n1846, ZN => n1871);
   U1294 : OAI21_X1 port map( B1 => n5477, B2 => n5863, A => n1872, ZN => n3748
                           );
   U1295 : NAND2_X1 port map( A1 => n346, A2 => n1846, ZN => n1872);
   U1296 : OAI21_X1 port map( B1 => n5474, B2 => n5863, A => n1873, ZN => n3747
                           );
   U1297 : NAND2_X1 port map( A1 => n347, A2 => n1846, ZN => n1873);
   U1298 : OAI21_X1 port map( B1 => n5471, B2 => n5864, A => n1874, ZN => n3746
                           );
   U1299 : NAND2_X1 port map( A1 => n348, A2 => n1846, ZN => n1874);
   U1300 : OAI21_X1 port map( B1 => n5468, B2 => n5864, A => n1875, ZN => n3745
                           );
   U1301 : NAND2_X1 port map( A1 => n349, A2 => n5864, ZN => n1875);
   U1302 : OAI21_X1 port map( B1 => n5465, B2 => n5864, A => n1876, ZN => n3744
                           );
   U1303 : NAND2_X1 port map( A1 => n350, A2 => n5863, ZN => n1876);
   U1304 : OAI21_X1 port map( B1 => n5462, B2 => n5864, A => n1877, ZN => n3743
                           );
   U1305 : NAND2_X1 port map( A1 => n351, A2 => n1846, ZN => n1877);
   U1306 : OAI21_X1 port map( B1 => n5459, B2 => n1846, A => n1878, ZN => n3742
                           );
   U1307 : NAND2_X1 port map( A1 => n352, A2 => n5863, ZN => n1878);
   U1308 : NAND2_X1 port map( A1 => n1777, A2 => n1658, ZN => n1846);
   U1309 : OAI21_X1 port map( B1 => n5552, B2 => n1879, A => n1880, ZN => n3741
                           );
   U1310 : NAND2_X1 port map( A1 => n353, A2 => n5858, ZN => n1880);
   U1311 : OAI21_X1 port map( B1 => n5549, B2 => n1879, A => n1881, ZN => n3740
                           );
   U1312 : NAND2_X1 port map( A1 => n354, A2 => n5858, ZN => n1881);
   U1313 : OAI21_X1 port map( B1 => n5546, B2 => n1879, A => n1882, ZN => n3739
                           );
   U1314 : NAND2_X1 port map( A1 => n355, A2 => n5858, ZN => n1882);
   U1315 : OAI21_X1 port map( B1 => n5543, B2 => n1879, A => n1883, ZN => n3738
                           );
   U1316 : NAND2_X1 port map( A1 => n356, A2 => n5858, ZN => n1883);
   U1317 : OAI21_X1 port map( B1 => n5540, B2 => n1879, A => n1884, ZN => n3737
                           );
   U1318 : NAND2_X1 port map( A1 => n357, A2 => n5854, ZN => n1884);
   U1319 : OAI21_X1 port map( B1 => n5537, B2 => n1879, A => n1885, ZN => n3736
                           );
   U1320 : NAND2_X1 port map( A1 => n358, A2 => n5854, ZN => n1885);
   U1321 : OAI21_X1 port map( B1 => n5534, B2 => n1879, A => n1886, ZN => n3735
                           );
   U1322 : NAND2_X1 port map( A1 => n359, A2 => n5854, ZN => n1886);
   U1323 : OAI21_X1 port map( B1 => n5531, B2 => n1879, A => n1887, ZN => n3734
                           );
   U1324 : NAND2_X1 port map( A1 => n360, A2 => n1879, ZN => n1887);
   U1325 : OAI21_X1 port map( B1 => n5528, B2 => n1879, A => n1888, ZN => n3733
                           );
   U1326 : NAND2_X1 port map( A1 => n361, A2 => n1879, ZN => n1888);
   U1327 : OAI21_X1 port map( B1 => n6081, B2 => n1879, A => n1889, ZN => n3732
                           );
   U1328 : NAND2_X1 port map( A1 => n362, A2 => n1879, ZN => n1889);
   U1329 : OAI21_X1 port map( B1 => n5522, B2 => n1879, A => n1890, ZN => n3731
                           );
   U1330 : NAND2_X1 port map( A1 => n363, A2 => n1879, ZN => n1890);
   U1331 : OAI21_X1 port map( B1 => n5519, B2 => n1879, A => n1891, ZN => n3730
                           );
   U1332 : NAND2_X1 port map( A1 => n364, A2 => n1879, ZN => n1891);
   U1333 : OAI21_X1 port map( B1 => n5516, B2 => n1879, A => n1892, ZN => n3729
                           );
   U1334 : NAND2_X1 port map( A1 => n365, A2 => n5858, ZN => n1892);
   U1335 : OAI21_X1 port map( B1 => n5513, B2 => n1879, A => n1893, ZN => n3728
                           );
   U1336 : NAND2_X1 port map( A1 => n366, A2 => n5854, ZN => n1893);
   U1337 : OAI21_X1 port map( B1 => n5509, B2 => n1879, A => n1894, ZN => n3727
                           );
   U1338 : NAND2_X1 port map( A1 => n367, A2 => n1879, ZN => n1894);
   U1339 : OAI21_X1 port map( B1 => n5506, B2 => n5858, A => n1895, ZN => n3726
                           );
   U1340 : NAND2_X1 port map( A1 => n368, A2 => n1879, ZN => n1895);
   U1341 : OAI21_X1 port map( B1 => n5504, B2 => n5854, A => n1896, ZN => n3725
                           );
   U1342 : NAND2_X1 port map( A1 => n369, A2 => n5854, ZN => n1896);
   U1343 : OAI21_X1 port map( B1 => n6073, B2 => n5858, A => n1897, ZN => n3724
                           );
   U1344 : NAND2_X1 port map( A1 => n370, A2 => n5854, ZN => n1897);
   U1345 : OAI21_X1 port map( B1 => n5498, B2 => n5854, A => n1898, ZN => n3723
                           );
   U1346 : NAND2_X1 port map( A1 => n371, A2 => n5854, ZN => n1898);
   U1347 : OAI21_X1 port map( B1 => n5495, B2 => n5858, A => n1899, ZN => n3722
                           );
   U1348 : NAND2_X1 port map( A1 => n372, A2 => n5854, ZN => n1899);
   U1349 : OAI21_X1 port map( B1 => n5492, B2 => n5854, A => n1900, ZN => n3721
                           );
   U1350 : NAND2_X1 port map( A1 => n373, A2 => n5854, ZN => n1900);
   U1351 : OAI21_X1 port map( B1 => n5489, B2 => n5858, A => n1901, ZN => n3720
                           );
   U1352 : NAND2_X1 port map( A1 => n374, A2 => n5854, ZN => n1901);
   U1353 : OAI21_X1 port map( B1 => n5486, B2 => n5854, A => n1902, ZN => n3719
                           );
   U1354 : NAND2_X1 port map( A1 => n375, A2 => n5854, ZN => n1902);
   U1355 : OAI21_X1 port map( B1 => n6067, B2 => n5858, A => n1903, ZN => n3718
                           );
   U1356 : NAND2_X1 port map( A1 => n376, A2 => n5854, ZN => n1903);
   U1357 : OAI21_X1 port map( B1 => n5480, B2 => n5854, A => n1904, ZN => n3717
                           );
   U1358 : NAND2_X1 port map( A1 => n377, A2 => n5858, ZN => n1904);
   U1359 : OAI21_X1 port map( B1 => n5477, B2 => n5858, A => n1905, ZN => n3716
                           );
   U1360 : NAND2_X1 port map( A1 => n378, A2 => n5858, ZN => n1905);
   U1361 : OAI21_X1 port map( B1 => n5474, B2 => n5854, A => n1906, ZN => n3715
                           );
   U1362 : NAND2_X1 port map( A1 => n379, A2 => n5858, ZN => n1906);
   U1363 : OAI21_X1 port map( B1 => n5471, B2 => n5858, A => n1907, ZN => n3714
                           );
   U1364 : NAND2_X1 port map( A1 => n380, A2 => n5858, ZN => n1907);
   U1365 : OAI21_X1 port map( B1 => n5468, B2 => n5858, A => n1908, ZN => n3713
                           );
   U1366 : NAND2_X1 port map( A1 => n381, A2 => n5854, ZN => n1908);
   U1367 : OAI21_X1 port map( B1 => n5465, B2 => n5858, A => n1909, ZN => n3712
                           );
   U1368 : NAND2_X1 port map( A1 => n382, A2 => n5854, ZN => n1909);
   U1369 : OAI21_X1 port map( B1 => n5462, B2 => n5858, A => n1910, ZN => n3711
                           );
   U1370 : NAND2_X1 port map( A1 => n383, A2 => n1879, ZN => n1910);
   U1371 : OAI21_X1 port map( B1 => n5459, B2 => n1879, A => n1911, ZN => n3710
                           );
   U1372 : NAND2_X1 port map( A1 => n384, A2 => n5858, ZN => n1911);
   U1373 : NAND2_X1 port map( A1 => n1777, A2 => n1624, ZN => n1879);
   U1374 : OAI21_X1 port map( B1 => n5552, B2 => n5850, A => n1913, ZN => n3709
                           );
   U1375 : NAND2_X1 port map( A1 => n641, A2 => n1912, ZN => n1913);
   U1376 : OAI21_X1 port map( B1 => n5549, B2 => n5850, A => n1914, ZN => n3708
                           );
   U1377 : NAND2_X1 port map( A1 => n642, A2 => n1912, ZN => n1914);
   U1378 : OAI21_X1 port map( B1 => n5546, B2 => n5850, A => n1915, ZN => n3707
                           );
   U1379 : NAND2_X1 port map( A1 => n643, A2 => n1912, ZN => n1915);
   U1380 : OAI21_X1 port map( B1 => n5543, B2 => n5851, A => n1916, ZN => n3706
                           );
   U1381 : NAND2_X1 port map( A1 => n644, A2 => n1912, ZN => n1916);
   U1382 : OAI21_X1 port map( B1 => n5540, B2 => n5850, A => n1917, ZN => n3705
                           );
   U1383 : NAND2_X1 port map( A1 => n645, A2 => n5851, ZN => n1917);
   U1384 : OAI21_X1 port map( B1 => n5537, B2 => n5850, A => n1918, ZN => n3704
                           );
   U1385 : NAND2_X1 port map( A1 => n646, A2 => n1912, ZN => n1918);
   U1386 : OAI21_X1 port map( B1 => n5534, B2 => n5850, A => n1919, ZN => n3703
                           );
   U1387 : NAND2_X1 port map( A1 => n647, A2 => n1912, ZN => n1919);
   U1388 : OAI21_X1 port map( B1 => n5531, B2 => n5850, A => n1920, ZN => n3702
                           );
   U1389 : NAND2_X1 port map( A1 => n648, A2 => n5850, ZN => n1920);
   U1390 : OAI21_X1 port map( B1 => n5528, B2 => n5850, A => n1921, ZN => n3701
                           );
   U1391 : NAND2_X1 port map( A1 => n649, A2 => n5851, ZN => n1921);
   U1392 : OAI21_X1 port map( B1 => n6081, B2 => n5850, A => n1922, ZN => n3700
                           );
   U1393 : NAND2_X1 port map( A1 => n650, A2 => n5850, ZN => n1922);
   U1394 : OAI21_X1 port map( B1 => n5522, B2 => n5850, A => n1923, ZN => n3699
                           );
   U1395 : NAND2_X1 port map( A1 => n651, A2 => n5851, ZN => n1923);
   U1396 : OAI21_X1 port map( B1 => n5519, B2 => n5850, A => n1924, ZN => n3698
                           );
   U1397 : NAND2_X1 port map( A1 => n652, A2 => n5850, ZN => n1924);
   U1398 : OAI21_X1 port map( B1 => n5516, B2 => n5850, A => n1925, ZN => n3697
                           );
   U1399 : NAND2_X1 port map( A1 => n653, A2 => n5851, ZN => n1925);
   U1400 : OAI21_X1 port map( B1 => n5513, B2 => n5850, A => n1926, ZN => n3696
                           );
   U1401 : NAND2_X1 port map( A1 => n654, A2 => n1912, ZN => n1926);
   U1402 : OAI21_X1 port map( B1 => n5509, B2 => n5850, A => n1927, ZN => n3695
                           );
   U1403 : NAND2_X1 port map( A1 => n655, A2 => n5850, ZN => n1927);
   U1404 : OAI21_X1 port map( B1 => n5506, B2 => n5851, A => n1928, ZN => n3694
                           );
   U1405 : NAND2_X1 port map( A1 => n656, A2 => n5850, ZN => n1928);
   U1406 : OAI21_X1 port map( B1 => n5504, B2 => n5851, A => n1929, ZN => n3693
                           );
   U1407 : NAND2_X1 port map( A1 => n657, A2 => n1912, ZN => n1929);
   U1408 : OAI21_X1 port map( B1 => n6073, B2 => n5851, A => n1930, ZN => n3692
                           );
   U1409 : NAND2_X1 port map( A1 => n658, A2 => n1912, ZN => n1930);
   U1410 : OAI21_X1 port map( B1 => n5498, B2 => n5851, A => n1931, ZN => n3691
                           );
   U1411 : NAND2_X1 port map( A1 => n659, A2 => n1912, ZN => n1931);
   U1412 : OAI21_X1 port map( B1 => n5495, B2 => n5851, A => n1932, ZN => n3690
                           );
   U1413 : NAND2_X1 port map( A1 => n660, A2 => n1912, ZN => n1932);
   U1414 : OAI21_X1 port map( B1 => n5492, B2 => n5851, A => n1933, ZN => n3689
                           );
   U1415 : NAND2_X1 port map( A1 => n661, A2 => n1912, ZN => n1933);
   U1416 : OAI21_X1 port map( B1 => n5489, B2 => n5851, A => n1934, ZN => n3688
                           );
   U1417 : NAND2_X1 port map( A1 => n662, A2 => n1912, ZN => n1934);
   U1418 : OAI21_X1 port map( B1 => n5486, B2 => n5851, A => n1935, ZN => n3687
                           );
   U1419 : NAND2_X1 port map( A1 => n663, A2 => n1912, ZN => n1935);
   U1420 : OAI21_X1 port map( B1 => n6067, B2 => n5851, A => n1936, ZN => n3686
                           );
   U1421 : NAND2_X1 port map( A1 => n664, A2 => n1912, ZN => n1936);
   U1422 : OAI21_X1 port map( B1 => n5480, B2 => n5851, A => n1937, ZN => n3685
                           );
   U1423 : NAND2_X1 port map( A1 => n665, A2 => n1912, ZN => n1937);
   U1424 : OAI21_X1 port map( B1 => n5477, B2 => n5851, A => n1938, ZN => n3684
                           );
   U1425 : NAND2_X1 port map( A1 => n666, A2 => n1912, ZN => n1938);
   U1426 : OAI21_X1 port map( B1 => n5474, B2 => n5851, A => n1939, ZN => n3683
                           );
   U1427 : NAND2_X1 port map( A1 => n667, A2 => n1912, ZN => n1939);
   U1428 : OAI21_X1 port map( B1 => n5471, B2 => n5850, A => n1940, ZN => n3682
                           );
   U1429 : NAND2_X1 port map( A1 => n668, A2 => n1912, ZN => n1940);
   U1430 : OAI21_X1 port map( B1 => n5468, B2 => n5851, A => n1941, ZN => n3681
                           );
   U1431 : NAND2_X1 port map( A1 => n669, A2 => n1912, ZN => n1941);
   U1432 : OAI21_X1 port map( B1 => n5465, B2 => n5850, A => n1942, ZN => n3680
                           );
   U1433 : NAND2_X1 port map( A1 => n670, A2 => n1912, ZN => n1942);
   U1434 : OAI21_X1 port map( B1 => n5462, B2 => n5851, A => n1943, ZN => n3679
                           );
   U1435 : NAND2_X1 port map( A1 => n671, A2 => n1912, ZN => n1943);
   U1436 : OAI21_X1 port map( B1 => n5459, B2 => n5851, A => n1944, ZN => n3678
                           );
   U1437 : NAND2_X1 port map( A1 => n672, A2 => n1912, ZN => n1944);
   U1438 : NAND2_X1 port map( A1 => n1777, A2 => n1590, ZN => n1912);
   U1439 : OAI21_X1 port map( B1 => n5552, B2 => n5846, A => n1946, ZN => n3677
                           );
   U1440 : NAND2_X1 port map( A1 => n481, A2 => n1945, ZN => n1946);
   U1441 : OAI21_X1 port map( B1 => n5549, B2 => n1945, A => n1947, ZN => n3676
                           );
   U1442 : NAND2_X1 port map( A1 => n482, A2 => n1945, ZN => n1947);
   U1443 : OAI21_X1 port map( B1 => n5546, B2 => n5845, A => n1948, ZN => n3675
                           );
   U1444 : NAND2_X1 port map( A1 => n483, A2 => n1945, ZN => n1948);
   U1445 : OAI21_X1 port map( B1 => n5543, B2 => n1945, A => n1949, ZN => n3674
                           );
   U1446 : NAND2_X1 port map( A1 => n484, A2 => n1945, ZN => n1949);
   U1447 : OAI21_X1 port map( B1 => n5540, B2 => n1945, A => n1950, ZN => n3673
                           );
   U1448 : NAND2_X1 port map( A1 => n485, A2 => n5846, ZN => n1950);
   U1449 : OAI21_X1 port map( B1 => n5537, B2 => n5846, A => n1951, ZN => n3672
                           );
   U1450 : NAND2_X1 port map( A1 => n486, A2 => n5846, ZN => n1951);
   U1451 : OAI21_X1 port map( B1 => n5534, B2 => n5845, A => n1952, ZN => n3671
                           );
   U1452 : NAND2_X1 port map( A1 => n487, A2 => n1945, ZN => n1952);
   U1453 : OAI21_X1 port map( B1 => n5531, B2 => n5846, A => n1953, ZN => n3670
                           );
   U1454 : NAND2_X1 port map( A1 => n488, A2 => n1945, ZN => n1953);
   U1455 : OAI21_X1 port map( B1 => n5528, B2 => n5845, A => n1954, ZN => n3669
                           );
   U1456 : NAND2_X1 port map( A1 => n489, A2 => n1945, ZN => n1954);
   U1457 : OAI21_X1 port map( B1 => n6081, B2 => n5846, A => n1955, ZN => n3668
                           );
   U1458 : NAND2_X1 port map( A1 => n490, A2 => n1945, ZN => n1955);
   U1459 : OAI21_X1 port map( B1 => n5522, B2 => n5845, A => n1956, ZN => n3667
                           );
   U1460 : NAND2_X1 port map( A1 => n491, A2 => n1945, ZN => n1956);
   U1461 : OAI21_X1 port map( B1 => n5519, B2 => n5846, A => n1957, ZN => n3666
                           );
   U1462 : NAND2_X1 port map( A1 => n492, A2 => n1945, ZN => n1957);
   U1463 : OAI21_X1 port map( B1 => n5516, B2 => n5845, A => n1958, ZN => n3665
                           );
   U1464 : NAND2_X1 port map( A1 => n493, A2 => n1945, ZN => n1958);
   U1465 : OAI21_X1 port map( B1 => n5513, B2 => n1945, A => n1959, ZN => n3664
                           );
   U1466 : NAND2_X1 port map( A1 => n494, A2 => n5846, ZN => n1959);
   U1467 : OAI21_X1 port map( B1 => n5509, B2 => n1945, A => n1960, ZN => n3663
                           );
   U1468 : NAND2_X1 port map( A1 => n495, A2 => n1945, ZN => n1960);
   U1469 : OAI21_X1 port map( B1 => n5506, B2 => n5845, A => n1961, ZN => n3662
                           );
   U1470 : NAND2_X1 port map( A1 => n496, A2 => n1945, ZN => n1961);
   U1471 : OAI21_X1 port map( B1 => n5504, B2 => n5845, A => n1962, ZN => n3661
                           );
   U1472 : NAND2_X1 port map( A1 => n497, A2 => n5845, ZN => n1962);
   U1473 : OAI21_X1 port map( B1 => n6073, B2 => n5845, A => n1963, ZN => n3660
                           );
   U1474 : NAND2_X1 port map( A1 => n498, A2 => n5846, ZN => n1963);
   U1475 : OAI21_X1 port map( B1 => n5498, B2 => n5845, A => n1964, ZN => n3659
                           );
   U1476 : NAND2_X1 port map( A1 => n499, A2 => n5846, ZN => n1964);
   U1477 : OAI21_X1 port map( B1 => n5495, B2 => n5845, A => n1965, ZN => n3658
                           );
   U1478 : NAND2_X1 port map( A1 => n500, A2 => n5846, ZN => n1965);
   U1479 : OAI21_X1 port map( B1 => n5492, B2 => n5845, A => n1966, ZN => n3657
                           );
   U1480 : NAND2_X1 port map( A1 => n501, A2 => n5846, ZN => n1966);
   U1481 : OAI21_X1 port map( B1 => n5489, B2 => n5845, A => n1967, ZN => n3656
                           );
   U1482 : NAND2_X1 port map( A1 => n502, A2 => n5846, ZN => n1967);
   U1483 : OAI21_X1 port map( B1 => n5486, B2 => n5845, A => n1968, ZN => n3655
                           );
   U1484 : NAND2_X1 port map( A1 => n503, A2 => n5846, ZN => n1968);
   U1485 : OAI21_X1 port map( B1 => n6067, B2 => n5845, A => n1969, ZN => n3654
                           );
   U1486 : NAND2_X1 port map( A1 => n504, A2 => n5846, ZN => n1969);
   U1487 : OAI21_X1 port map( B1 => n5480, B2 => n5845, A => n1970, ZN => n3653
                           );
   U1488 : NAND2_X1 port map( A1 => n505, A2 => n1945, ZN => n1970);
   U1489 : OAI21_X1 port map( B1 => n5477, B2 => n5845, A => n1971, ZN => n3652
                           );
   U1490 : NAND2_X1 port map( A1 => n506, A2 => n1945, ZN => n1971);
   U1491 : OAI21_X1 port map( B1 => n5474, B2 => n5845, A => n1972, ZN => n3651
                           );
   U1492 : NAND2_X1 port map( A1 => n507, A2 => n1945, ZN => n1972);
   U1493 : OAI21_X1 port map( B1 => n5471, B2 => n5846, A => n1973, ZN => n3650
                           );
   U1494 : NAND2_X1 port map( A1 => n508, A2 => n1945, ZN => n1973);
   U1495 : OAI21_X1 port map( B1 => n5468, B2 => n5846, A => n1974, ZN => n3649
                           );
   U1496 : NAND2_X1 port map( A1 => n509, A2 => n5846, ZN => n1974);
   U1497 : OAI21_X1 port map( B1 => n5465, B2 => n5846, A => n1975, ZN => n3648
                           );
   U1498 : NAND2_X1 port map( A1 => n510, A2 => n5845, ZN => n1975);
   U1499 : OAI21_X1 port map( B1 => n5462, B2 => n5846, A => n1976, ZN => n3647
                           );
   U1500 : NAND2_X1 port map( A1 => n511, A2 => n1945, ZN => n1976);
   U1501 : OAI21_X1 port map( B1 => n5459, B2 => n1945, A => n1977, ZN => n3646
                           );
   U1502 : NAND2_X1 port map( A1 => n512, A2 => n5845, ZN => n1977);
   U1503 : NAND2_X1 port map( A1 => n1777, A2 => n1555, ZN => n1945);
   U1504 : OAI21_X1 port map( B1 => n5552, B2 => n5840, A => n1979, ZN => n3645
                           );
   U1505 : NAND2_X1 port map( A1 => n513, A2 => n1978, ZN => n1979);
   U1506 : OAI21_X1 port map( B1 => n5549, B2 => n1978, A => n1980, ZN => n3644
                           );
   U1507 : NAND2_X1 port map( A1 => n514, A2 => n1978, ZN => n1980);
   U1508 : OAI21_X1 port map( B1 => n5546, B2 => n5839, A => n1981, ZN => n3643
                           );
   U1509 : NAND2_X1 port map( A1 => n515, A2 => n1978, ZN => n1981);
   U1510 : OAI21_X1 port map( B1 => n5543, B2 => n1978, A => n1982, ZN => n3642
                           );
   U1511 : NAND2_X1 port map( A1 => n516, A2 => n1978, ZN => n1982);
   U1512 : OAI21_X1 port map( B1 => n5540, B2 => n1978, A => n1983, ZN => n3641
                           );
   U1513 : NAND2_X1 port map( A1 => n517, A2 => n5840, ZN => n1983);
   U1514 : OAI21_X1 port map( B1 => n5537, B2 => n5840, A => n1984, ZN => n3640
                           );
   U1515 : NAND2_X1 port map( A1 => n518, A2 => n5840, ZN => n1984);
   U1516 : OAI21_X1 port map( B1 => n5534, B2 => n5839, A => n1985, ZN => n3639
                           );
   U1517 : NAND2_X1 port map( A1 => n519, A2 => n1978, ZN => n1985);
   U1518 : OAI21_X1 port map( B1 => n5531, B2 => n5840, A => n1986, ZN => n3638
                           );
   U1519 : NAND2_X1 port map( A1 => n520, A2 => n1978, ZN => n1986);
   U1520 : OAI21_X1 port map( B1 => n5528, B2 => n5839, A => n1987, ZN => n3637
                           );
   U1521 : NAND2_X1 port map( A1 => n521, A2 => n1978, ZN => n1987);
   U1522 : OAI21_X1 port map( B1 => n6081, B2 => n5840, A => n1988, ZN => n3636
                           );
   U1523 : NAND2_X1 port map( A1 => n522, A2 => n1978, ZN => n1988);
   U1524 : OAI21_X1 port map( B1 => n5522, B2 => n5839, A => n1989, ZN => n3635
                           );
   U1525 : NAND2_X1 port map( A1 => n523, A2 => n1978, ZN => n1989);
   U1526 : OAI21_X1 port map( B1 => n5519, B2 => n5840, A => n1990, ZN => n3634
                           );
   U1527 : NAND2_X1 port map( A1 => n524, A2 => n1978, ZN => n1990);
   U1528 : OAI21_X1 port map( B1 => n5516, B2 => n5839, A => n1991, ZN => n3633
                           );
   U1529 : NAND2_X1 port map( A1 => n525, A2 => n1978, ZN => n1991);
   U1530 : OAI21_X1 port map( B1 => n5513, B2 => n1978, A => n1992, ZN => n3632
                           );
   U1531 : NAND2_X1 port map( A1 => n526, A2 => n5840, ZN => n1992);
   U1532 : OAI21_X1 port map( B1 => n5509, B2 => n1978, A => n1993, ZN => n3631
                           );
   U1533 : NAND2_X1 port map( A1 => n527, A2 => n1978, ZN => n1993);
   U1534 : OAI21_X1 port map( B1 => n5506, B2 => n5839, A => n1994, ZN => n3630
                           );
   U1535 : NAND2_X1 port map( A1 => n528, A2 => n1978, ZN => n1994);
   U1536 : OAI21_X1 port map( B1 => n5504, B2 => n5839, A => n1995, ZN => n3629
                           );
   U1537 : NAND2_X1 port map( A1 => n529, A2 => n5839, ZN => n1995);
   U1538 : OAI21_X1 port map( B1 => n6073, B2 => n5839, A => n1996, ZN => n3628
                           );
   U1539 : NAND2_X1 port map( A1 => n530, A2 => n5840, ZN => n1996);
   U1540 : OAI21_X1 port map( B1 => n5498, B2 => n5839, A => n1997, ZN => n3627
                           );
   U1541 : NAND2_X1 port map( A1 => n531, A2 => n5840, ZN => n1997);
   U1542 : OAI21_X1 port map( B1 => n5495, B2 => n5839, A => n1998, ZN => n3626
                           );
   U1543 : NAND2_X1 port map( A1 => n532, A2 => n5840, ZN => n1998);
   U1544 : OAI21_X1 port map( B1 => n5492, B2 => n5839, A => n1999, ZN => n3625
                           );
   U1545 : NAND2_X1 port map( A1 => n533, A2 => n5840, ZN => n1999);
   U1546 : OAI21_X1 port map( B1 => n5489, B2 => n5839, A => n2000, ZN => n3624
                           );
   U1547 : NAND2_X1 port map( A1 => n534, A2 => n5840, ZN => n2000);
   U1548 : OAI21_X1 port map( B1 => n5486, B2 => n5839, A => n2001, ZN => n3623
                           );
   U1549 : NAND2_X1 port map( A1 => n535, A2 => n5840, ZN => n2001);
   U1550 : OAI21_X1 port map( B1 => n6067, B2 => n5839, A => n2002, ZN => n3622
                           );
   U1551 : NAND2_X1 port map( A1 => n536, A2 => n5840, ZN => n2002);
   U1552 : OAI21_X1 port map( B1 => n5480, B2 => n5839, A => n2003, ZN => n3621
                           );
   U1553 : NAND2_X1 port map( A1 => n537, A2 => n1978, ZN => n2003);
   U1554 : OAI21_X1 port map( B1 => n5477, B2 => n5839, A => n2004, ZN => n3620
                           );
   U1555 : NAND2_X1 port map( A1 => n538, A2 => n1978, ZN => n2004);
   U1556 : OAI21_X1 port map( B1 => n5474, B2 => n5839, A => n2005, ZN => n3619
                           );
   U1557 : NAND2_X1 port map( A1 => n539, A2 => n1978, ZN => n2005);
   U1558 : OAI21_X1 port map( B1 => n5471, B2 => n5840, A => n2006, ZN => n3618
                           );
   U1559 : NAND2_X1 port map( A1 => n540, A2 => n1978, ZN => n2006);
   U1560 : OAI21_X1 port map( B1 => n5468, B2 => n5840, A => n2007, ZN => n3617
                           );
   U1561 : NAND2_X1 port map( A1 => n541, A2 => n5840, ZN => n2007);
   U1562 : OAI21_X1 port map( B1 => n5465, B2 => n5840, A => n2008, ZN => n3616
                           );
   U1563 : NAND2_X1 port map( A1 => n542, A2 => n5839, ZN => n2008);
   U1564 : OAI21_X1 port map( B1 => n5462, B2 => n5840, A => n2009, ZN => n3615
                           );
   U1565 : NAND2_X1 port map( A1 => n543, A2 => n1978, ZN => n2009);
   U1566 : OAI21_X1 port map( B1 => n5459, B2 => n1978, A => n2010, ZN => n3614
                           );
   U1567 : NAND2_X1 port map( A1 => n544, A2 => n5839, ZN => n2010);
   U1568 : NAND2_X1 port map( A1 => n1692, A2 => n1521, ZN => n1978);
   U1569 : OAI21_X1 port map( B1 => n5552, B2 => n5829, A => n2012, ZN => n3613
                           );
   U1570 : NAND2_X1 port map( A1 => n705, A2 => n5829, ZN => n2012);
   U1571 : OAI21_X1 port map( B1 => n5549, B2 => n5831, A => n2013, ZN => n3612
                           );
   U1572 : NAND2_X1 port map( A1 => n706, A2 => n5829, ZN => n2013);
   U1573 : OAI21_X1 port map( B1 => n5546, B2 => n2011, A => n2014, ZN => n3611
                           );
   U1574 : NAND2_X1 port map( A1 => n707, A2 => n5829, ZN => n2014);
   U1575 : OAI21_X1 port map( B1 => n5543, B2 => n5831, A => n2015, ZN => n3610
                           );
   U1576 : NAND2_X1 port map( A1 => n708, A2 => n5829, ZN => n2015);
   U1577 : OAI21_X1 port map( B1 => n5540, B2 => n5831, A => n2016, ZN => n3609
                           );
   U1578 : NAND2_X1 port map( A1 => n709, A2 => n5831, ZN => n2016);
   U1579 : OAI21_X1 port map( B1 => n5537, B2 => n2011, A => n2017, ZN => n3608
                           );
   U1580 : NAND2_X1 port map( A1 => n710, A2 => n5831, ZN => n2017);
   U1581 : OAI21_X1 port map( B1 => n5534, B2 => n2011, A => n2018, ZN => n3607
                           );
   U1582 : NAND2_X1 port map( A1 => n711, A2 => n5829, ZN => n2018);
   U1583 : OAI21_X1 port map( B1 => n5531, B2 => n2011, A => n2019, ZN => n3606
                           );
   U1584 : NAND2_X1 port map( A1 => n712, A2 => n5831, ZN => n2019);
   U1585 : OAI21_X1 port map( B1 => n5528, B2 => n2011, A => n2020, ZN => n3605
                           );
   U1586 : NAND2_X1 port map( A1 => n713, A2 => n5831, ZN => n2020);
   U1587 : OAI21_X1 port map( B1 => n6081, B2 => n2011, A => n2021, ZN => n3604
                           );
   U1588 : NAND2_X1 port map( A1 => n714, A2 => n5831, ZN => n2021);
   U1589 : OAI21_X1 port map( B1 => n5522, B2 => n2011, A => n2022, ZN => n3603
                           );
   U1590 : NAND2_X1 port map( A1 => n715, A2 => n5831, ZN => n2022);
   U1591 : OAI21_X1 port map( B1 => n5519, B2 => n2011, A => n2023, ZN => n3602
                           );
   U1592 : NAND2_X1 port map( A1 => n716, A2 => n5831, ZN => n2023);
   U1593 : OAI21_X1 port map( B1 => n5516, B2 => n2011, A => n2024, ZN => n3601
                           );
   U1594 : NAND2_X1 port map( A1 => n717, A2 => n5831, ZN => n2024);
   U1595 : OAI21_X1 port map( B1 => n5513, B2 => n2011, A => n2025, ZN => n3600
                           );
   U1596 : NAND2_X1 port map( A1 => n718, A2 => n5831, ZN => n2025);
   U1597 : OAI21_X1 port map( B1 => n5509, B2 => n2011, A => n2026, ZN => n3599
                           );
   U1598 : NAND2_X1 port map( A1 => n719, A2 => n5831, ZN => n2026);
   U1599 : OAI21_X1 port map( B1 => n5506, B2 => n2011, A => n2027, ZN => n3598
                           );
   U1600 : NAND2_X1 port map( A1 => n720, A2 => n5831, ZN => n2027);
   U1601 : OAI21_X1 port map( B1 => n5504, B2 => n2011, A => n2028, ZN => n3597
                           );
   U1602 : NAND2_X1 port map( A1 => n721, A2 => n5829, ZN => n2028);
   U1603 : OAI21_X1 port map( B1 => n6073, B2 => n2011, A => n2029, ZN => n3596
                           );
   U1604 : NAND2_X1 port map( A1 => n722, A2 => n5831, ZN => n2029);
   U1605 : OAI21_X1 port map( B1 => n5498, B2 => n2011, A => n2030, ZN => n3595
                           );
   U1606 : NAND2_X1 port map( A1 => n723, A2 => n5829, ZN => n2030);
   U1607 : OAI21_X1 port map( B1 => n5495, B2 => n2011, A => n2031, ZN => n3594
                           );
   U1608 : NAND2_X1 port map( A1 => n724, A2 => n5831, ZN => n2031);
   U1609 : OAI21_X1 port map( B1 => n5492, B2 => n2011, A => n2032, ZN => n3593
                           );
   U1610 : NAND2_X1 port map( A1 => n725, A2 => n5829, ZN => n2032);
   U1611 : OAI21_X1 port map( B1 => n5489, B2 => n2011, A => n2033, ZN => n3592
                           );
   U1612 : NAND2_X1 port map( A1 => n726, A2 => n5831, ZN => n2033);
   U1613 : OAI21_X1 port map( B1 => n5486, B2 => n2011, A => n2034, ZN => n3591
                           );
   U1614 : NAND2_X1 port map( A1 => n727, A2 => n5829, ZN => n2034);
   U1615 : OAI21_X1 port map( B1 => n6067, B2 => n2011, A => n2035, ZN => n3590
                           );
   U1616 : NAND2_X1 port map( A1 => n728, A2 => n5831, ZN => n2035);
   U1617 : OAI21_X1 port map( B1 => n5480, B2 => n5831, A => n2036, ZN => n3589
                           );
   U1618 : NAND2_X1 port map( A1 => n729, A2 => n5829, ZN => n2036);
   U1619 : OAI21_X1 port map( B1 => n5477, B2 => n2011, A => n2037, ZN => n3588
                           );
   U1620 : NAND2_X1 port map( A1 => n730, A2 => n5829, ZN => n2037);
   U1621 : OAI21_X1 port map( B1 => n5474, B2 => n2011, A => n2038, ZN => n3587
                           );
   U1622 : NAND2_X1 port map( A1 => n731, A2 => n5829, ZN => n2038);
   U1623 : OAI21_X1 port map( B1 => n5471, B2 => n2011, A => n2039, ZN => n3586
                           );
   U1624 : NAND2_X1 port map( A1 => n732, A2 => n5829, ZN => n2039);
   U1625 : OAI21_X1 port map( B1 => n5468, B2 => n2011, A => n2040, ZN => n3585
                           );
   U1626 : NAND2_X1 port map( A1 => n733, A2 => n5829, ZN => n2040);
   U1627 : OAI21_X1 port map( B1 => n5465, B2 => n5829, A => n2041, ZN => n3584
                           );
   U1628 : NAND2_X1 port map( A1 => n734, A2 => n5829, ZN => n2041);
   U1629 : OAI21_X1 port map( B1 => n5462, B2 => n5829, A => n2042, ZN => n3583
                           );
   U1630 : NAND2_X1 port map( A1 => n735, A2 => n5829, ZN => n2042);
   U1631 : OAI21_X1 port map( B1 => n5459, B2 => n5831, A => n2043, ZN => n3582
                           );
   U1632 : NAND2_X1 port map( A1 => n736, A2 => n5829, ZN => n2043);
   U1633 : NAND2_X1 port map( A1 => n1812, A2 => n1692, ZN => n2011);
   U1634 : OAI21_X1 port map( B1 => n5552, B2 => n5828, A => n2045, ZN => n3581
                           );
   U1635 : NAND2_X1 port map( A1 => n2044, A2 => n6635, ZN => n2045);
   U1636 : OAI21_X1 port map( B1 => n5549, B2 => n2044, A => n2046, ZN => n3580
                           );
   U1637 : NAND2_X1 port map( A1 => n2044, A2 => n6634, ZN => n2046);
   U1638 : OAI21_X1 port map( B1 => n5546, B2 => n5827, A => n2047, ZN => n3579
                           );
   U1639 : NAND2_X1 port map( A1 => n2044, A2 => n6633, ZN => n2047);
   U1640 : OAI21_X1 port map( B1 => n5543, B2 => n2044, A => n2048, ZN => n3578
                           );
   U1641 : NAND2_X1 port map( A1 => n2044, A2 => n6632, ZN => n2048);
   U1642 : OAI21_X1 port map( B1 => n5540, B2 => n2044, A => n2049, ZN => n3577
                           );
   U1643 : NAND2_X1 port map( A1 => n5828, A2 => n6631, ZN => n2049);
   U1644 : OAI21_X1 port map( B1 => n5537, B2 => n5828, A => n2050, ZN => n3576
                           );
   U1645 : NAND2_X1 port map( A1 => n2044, A2 => n6630, ZN => n2050);
   U1646 : OAI21_X1 port map( B1 => n5534, B2 => n5827, A => n2051, ZN => n3575
                           );
   U1647 : NAND2_X1 port map( A1 => n2044, A2 => n6629, ZN => n2051);
   U1648 : OAI21_X1 port map( B1 => n5531, B2 => n5828, A => n2052, ZN => n3574
                           );
   U1649 : NAND2_X1 port map( A1 => n2044, A2 => n6628, ZN => n2052);
   U1650 : OAI21_X1 port map( B1 => n5528, B2 => n5827, A => n2053, ZN => n3573
                           );
   U1651 : NAND2_X1 port map( A1 => n2044, A2 => n6627, ZN => n2053);
   U1652 : OAI21_X1 port map( B1 => n6081, B2 => n5828, A => n2054, ZN => n3572
                           );
   U1653 : NAND2_X1 port map( A1 => n2044, A2 => n6626, ZN => n2054);
   U1654 : OAI21_X1 port map( B1 => n5522, B2 => n5827, A => n2055, ZN => n3571
                           );
   U1655 : NAND2_X1 port map( A1 => n2044, A2 => n6625, ZN => n2055);
   U1656 : OAI21_X1 port map( B1 => n5519, B2 => n5828, A => n2056, ZN => n3570
                           );
   U1657 : NAND2_X1 port map( A1 => n2044, A2 => n6624, ZN => n2056);
   U1658 : OAI21_X1 port map( B1 => n5516, B2 => n5827, A => n2057, ZN => n3569
                           );
   U1659 : NAND2_X1 port map( A1 => n2044, A2 => n6623, ZN => n2057);
   U1660 : OAI21_X1 port map( B1 => n5513, B2 => n5828, A => n2058, ZN => n3568
                           );
   U1661 : NAND2_X1 port map( A1 => n2044, A2 => n6622, ZN => n2058);
   U1662 : OAI21_X1 port map( B1 => n5509, B2 => n2044, A => n2059, ZN => n3567
                           );
   U1663 : NAND2_X1 port map( A1 => n5827, A2 => n6621, ZN => n2059);
   U1664 : OAI21_X1 port map( B1 => n5506, B2 => n5827, A => n2060, ZN => n3566
                           );
   U1665 : NAND2_X1 port map( A1 => n5827, A2 => n6620, ZN => n2060);
   U1666 : OAI21_X1 port map( B1 => n5504, B2 => n5827, A => n2061, ZN => n3565
                           );
   U1667 : NAND2_X1 port map( A1 => n5827, A2 => n6619, ZN => n2061);
   U1668 : OAI21_X1 port map( B1 => n6073, B2 => n5827, A => n2062, ZN => n3564
                           );
   U1669 : NAND2_X1 port map( A1 => n5828, A2 => n6618, ZN => n2062);
   U1670 : OAI21_X1 port map( B1 => n5498, B2 => n5827, A => n2063, ZN => n3563
                           );
   U1671 : NAND2_X1 port map( A1 => n5828, A2 => n6617, ZN => n2063);
   U1672 : OAI21_X1 port map( B1 => n5495, B2 => n5827, A => n2064, ZN => n3562
                           );
   U1673 : NAND2_X1 port map( A1 => n5828, A2 => n6616, ZN => n2064);
   U1674 : OAI21_X1 port map( B1 => n5492, B2 => n5827, A => n2065, ZN => n3561
                           );
   U1675 : NAND2_X1 port map( A1 => n5828, A2 => n6615, ZN => n2065);
   U1676 : OAI21_X1 port map( B1 => n5489, B2 => n5827, A => n2066, ZN => n3560
                           );
   U1677 : NAND2_X1 port map( A1 => n5828, A2 => n6614, ZN => n2066);
   U1678 : OAI21_X1 port map( B1 => n5486, B2 => n5827, A => n2067, ZN => n3559
                           );
   U1679 : NAND2_X1 port map( A1 => n5828, A2 => n6613, ZN => n2067);
   U1680 : OAI21_X1 port map( B1 => n6067, B2 => n5827, A => n2068, ZN => n3558
                           );
   U1681 : NAND2_X1 port map( A1 => n5828, A2 => n6612, ZN => n2068);
   U1682 : OAI21_X1 port map( B1 => n5480, B2 => n5827, A => n2069, ZN => n3557
                           );
   U1683 : NAND2_X1 port map( A1 => n5828, A2 => n6611, ZN => n2069);
   U1684 : OAI21_X1 port map( B1 => n5477, B2 => n5827, A => n2070, ZN => n3556
                           );
   U1685 : NAND2_X1 port map( A1 => n2044, A2 => n6610, ZN => n2070);
   U1686 : OAI21_X1 port map( B1 => n5474, B2 => n5827, A => n2071, ZN => n3555
                           );
   U1687 : NAND2_X1 port map( A1 => n5828, A2 => n6609, ZN => n2071);
   U1688 : OAI21_X1 port map( B1 => n5471, B2 => n5828, A => n2072, ZN => n3554
                           );
   U1689 : NAND2_X1 port map( A1 => n2044, A2 => n6608, ZN => n2072);
   U1690 : OAI21_X1 port map( B1 => n5468, B2 => n5828, A => n2073, ZN => n3553
                           );
   U1691 : NAND2_X1 port map( A1 => n2044, A2 => n6607, ZN => n2073);
   U1692 : OAI21_X1 port map( B1 => n5465, B2 => n5828, A => n2074, ZN => n3552
                           );
   U1693 : NAND2_X1 port map( A1 => n2044, A2 => n6606, ZN => n2074);
   U1694 : OAI21_X1 port map( B1 => n5462, B2 => n5828, A => n2075, ZN => n3551
                           );
   U1695 : NAND2_X1 port map( A1 => n2044, A2 => n6605, ZN => n2075);
   U1696 : OAI21_X1 port map( B1 => n5459, B2 => n2044, A => n2076, ZN => n3550
                           );
   U1697 : NAND2_X1 port map( A1 => n2044, A2 => n6604, ZN => n2076);
   U1698 : NAND2_X1 port map( A1 => n1778, A2 => n1692, ZN => n2044);
   U1699 : OAI21_X1 port map( B1 => n5552, B2 => n2077, A => n2078, ZN => n3549
                           );
   U1700 : NAND2_X1 port map( A1 => n673, A2 => n5822, ZN => n2078);
   U1701 : OAI21_X1 port map( B1 => n5549, B2 => n2077, A => n2079, ZN => n3548
                           );
   U1702 : NAND2_X1 port map( A1 => n674, A2 => n5822, ZN => n2079);
   U1703 : OAI21_X1 port map( B1 => n5546, B2 => n2077, A => n2080, ZN => n3547
                           );
   U1704 : NAND2_X1 port map( A1 => n675, A2 => n5822, ZN => n2080);
   U1705 : OAI21_X1 port map( B1 => n5543, B2 => n2077, A => n2081, ZN => n3546
                           );
   U1706 : NAND2_X1 port map( A1 => n676, A2 => n5822, ZN => n2081);
   U1707 : OAI21_X1 port map( B1 => n5540, B2 => n2077, A => n2082, ZN => n3545
                           );
   U1708 : NAND2_X1 port map( A1 => n677, A2 => n5818, ZN => n2082);
   U1709 : OAI21_X1 port map( B1 => n5537, B2 => n2077, A => n2083, ZN => n3544
                           );
   U1710 : NAND2_X1 port map( A1 => n678, A2 => n5818, ZN => n2083);
   U1711 : OAI21_X1 port map( B1 => n5534, B2 => n2077, A => n2084, ZN => n3543
                           );
   U1712 : NAND2_X1 port map( A1 => n679, A2 => n5818, ZN => n2084);
   U1713 : OAI21_X1 port map( B1 => n5531, B2 => n2077, A => n2085, ZN => n3542
                           );
   U1714 : NAND2_X1 port map( A1 => n680, A2 => n2077, ZN => n2085);
   U1715 : OAI21_X1 port map( B1 => n5528, B2 => n2077, A => n2086, ZN => n3541
                           );
   U1716 : NAND2_X1 port map( A1 => n681, A2 => n2077, ZN => n2086);
   U1717 : OAI21_X1 port map( B1 => n6081, B2 => n2077, A => n2087, ZN => n3540
                           );
   U1718 : NAND2_X1 port map( A1 => n682, A2 => n2077, ZN => n2087);
   U1719 : OAI21_X1 port map( B1 => n5522, B2 => n2077, A => n2088, ZN => n3539
                           );
   U1720 : NAND2_X1 port map( A1 => n683, A2 => n2077, ZN => n2088);
   U1721 : OAI21_X1 port map( B1 => n5519, B2 => n2077, A => n2089, ZN => n3538
                           );
   U1722 : NAND2_X1 port map( A1 => n684, A2 => n2077, ZN => n2089);
   U1723 : OAI21_X1 port map( B1 => n5516, B2 => n2077, A => n2090, ZN => n3537
                           );
   U1724 : NAND2_X1 port map( A1 => n685, A2 => n2077, ZN => n2090);
   U1725 : OAI21_X1 port map( B1 => n5513, B2 => n2077, A => n2091, ZN => n3536
                           );
   U1726 : NAND2_X1 port map( A1 => n686, A2 => n5818, ZN => n2091);
   U1727 : OAI21_X1 port map( B1 => n5509, B2 => n2077, A => n2092, ZN => n3535
                           );
   U1728 : NAND2_X1 port map( A1 => n687, A2 => n5822, ZN => n2092);
   U1729 : OAI21_X1 port map( B1 => n5506, B2 => n5822, A => n2093, ZN => n3534
                           );
   U1730 : NAND2_X1 port map( A1 => n688, A2 => n2077, ZN => n2093);
   U1731 : OAI21_X1 port map( B1 => n5504, B2 => n5818, A => n2094, ZN => n3533
                           );
   U1732 : NAND2_X1 port map( A1 => n689, A2 => n5818, ZN => n2094);
   U1733 : OAI21_X1 port map( B1 => n6073, B2 => n5822, A => n2095, ZN => n3532
                           );
   U1734 : NAND2_X1 port map( A1 => n690, A2 => n5818, ZN => n2095);
   U1735 : OAI21_X1 port map( B1 => n5498, B2 => n5818, A => n2096, ZN => n3531
                           );
   U1736 : NAND2_X1 port map( A1 => n691, A2 => n5818, ZN => n2096);
   U1737 : OAI21_X1 port map( B1 => n5495, B2 => n5822, A => n2097, ZN => n3530
                           );
   U1738 : NAND2_X1 port map( A1 => n692, A2 => n5818, ZN => n2097);
   U1739 : OAI21_X1 port map( B1 => n5492, B2 => n5818, A => n2098, ZN => n3529
                           );
   U1740 : NAND2_X1 port map( A1 => n693, A2 => n5818, ZN => n2098);
   U1741 : OAI21_X1 port map( B1 => n5489, B2 => n5822, A => n2099, ZN => n3528
                           );
   U1742 : NAND2_X1 port map( A1 => n694, A2 => n5818, ZN => n2099);
   U1743 : OAI21_X1 port map( B1 => n5486, B2 => n5818, A => n2100, ZN => n3527
                           );
   U1744 : NAND2_X1 port map( A1 => n695, A2 => n5818, ZN => n2100);
   U1745 : OAI21_X1 port map( B1 => n6067, B2 => n5822, A => n2101, ZN => n3526
                           );
   U1746 : NAND2_X1 port map( A1 => n696, A2 => n5818, ZN => n2101);
   U1747 : OAI21_X1 port map( B1 => n5480, B2 => n5818, A => n2102, ZN => n3525
                           );
   U1748 : NAND2_X1 port map( A1 => n697, A2 => n5822, ZN => n2102);
   U1749 : OAI21_X1 port map( B1 => n5477, B2 => n5822, A => n2103, ZN => n3524
                           );
   U1750 : NAND2_X1 port map( A1 => n698, A2 => n5822, ZN => n2103);
   U1751 : OAI21_X1 port map( B1 => n5474, B2 => n5818, A => n2104, ZN => n3523
                           );
   U1752 : NAND2_X1 port map( A1 => n699, A2 => n5822, ZN => n2104);
   U1753 : OAI21_X1 port map( B1 => n5471, B2 => n5822, A => n2105, ZN => n3522
                           );
   U1754 : NAND2_X1 port map( A1 => n700, A2 => n5822, ZN => n2105);
   U1755 : OAI21_X1 port map( B1 => n5468, B2 => n5822, A => n2106, ZN => n3521
                           );
   U1756 : NAND2_X1 port map( A1 => n701, A2 => n5818, ZN => n2106);
   U1757 : OAI21_X1 port map( B1 => n5465, B2 => n5822, A => n2107, ZN => n3520
                           );
   U1758 : NAND2_X1 port map( A1 => n702, A2 => n5818, ZN => n2107);
   U1759 : OAI21_X1 port map( B1 => n5462, B2 => n5822, A => n2108, ZN => n3519
                           );
   U1760 : NAND2_X1 port map( A1 => n703, A2 => n2077, ZN => n2108);
   U1761 : OAI21_X1 port map( B1 => n5459, B2 => n2077, A => n2109, ZN => n3518
                           );
   U1762 : NAND2_X1 port map( A1 => n704, A2 => n5822, ZN => n2109);
   U1763 : NAND2_X1 port map( A1 => n2110, A2 => n1692, ZN => n2077);
   U1764 : OAI21_X1 port map( B1 => n5552, B2 => n2111, A => n2112, ZN => n3517
                           );
   U1765 : NAND2_X1 port map( A1 => n5816, A2 => n6827, ZN => n2112);
   U1766 : OAI21_X1 port map( B1 => n5549, B2 => n2111, A => n2113, ZN => n3516
                           );
   U1767 : NAND2_X1 port map( A1 => n5816, A2 => n6826, ZN => n2113);
   U1768 : OAI21_X1 port map( B1 => n5546, B2 => n2111, A => n2114, ZN => n3515
                           );
   U1769 : NAND2_X1 port map( A1 => n5816, A2 => n6825, ZN => n2114);
   U1770 : OAI21_X1 port map( B1 => n5543, B2 => n2111, A => n2115, ZN => n3514
                           );
   U1771 : NAND2_X1 port map( A1 => n5816, A2 => n6824, ZN => n2115);
   U1772 : OAI21_X1 port map( B1 => n5540, B2 => n2111, A => n2116, ZN => n3513
                           );
   U1773 : NAND2_X1 port map( A1 => n5812, A2 => n6823, ZN => n2116);
   U1774 : OAI21_X1 port map( B1 => n5537, B2 => n2111, A => n2117, ZN => n3512
                           );
   U1775 : NAND2_X1 port map( A1 => n5812, A2 => n6822, ZN => n2117);
   U1776 : OAI21_X1 port map( B1 => n5534, B2 => n2111, A => n2118, ZN => n3511
                           );
   U1777 : NAND2_X1 port map( A1 => n5812, A2 => n6821, ZN => n2118);
   U1778 : OAI21_X1 port map( B1 => n5531, B2 => n2111, A => n2119, ZN => n3510
                           );
   U1779 : NAND2_X1 port map( A1 => n2111, A2 => n6820, ZN => n2119);
   U1780 : OAI21_X1 port map( B1 => n5528, B2 => n2111, A => n2120, ZN => n3509
                           );
   U1781 : NAND2_X1 port map( A1 => n2111, A2 => n6819, ZN => n2120);
   U1782 : OAI21_X1 port map( B1 => n6081, B2 => n2111, A => n2121, ZN => n3508
                           );
   U1783 : NAND2_X1 port map( A1 => n2111, A2 => n6818, ZN => n2121);
   U1784 : OAI21_X1 port map( B1 => n5522, B2 => n2111, A => n2122, ZN => n3507
                           );
   U1785 : NAND2_X1 port map( A1 => n2111, A2 => n6817, ZN => n2122);
   U1786 : OAI21_X1 port map( B1 => n5519, B2 => n2111, A => n2123, ZN => n3506
                           );
   U1787 : NAND2_X1 port map( A1 => n5812, A2 => n6816, ZN => n2123);
   U1788 : OAI21_X1 port map( B1 => n5516, B2 => n2111, A => n2124, ZN => n3505
                           );
   U1789 : NAND2_X1 port map( A1 => n5816, A2 => n6815, ZN => n2124);
   U1790 : OAI21_X1 port map( B1 => n5513, B2 => n2111, A => n2125, ZN => n3504
                           );
   U1791 : NAND2_X1 port map( A1 => n5812, A2 => n6814, ZN => n2125);
   U1792 : OAI21_X1 port map( B1 => n5509, B2 => n2111, A => n2126, ZN => n3503
                           );
   U1793 : NAND2_X1 port map( A1 => n2111, A2 => n6813, ZN => n2126);
   U1794 : OAI21_X1 port map( B1 => n5506, B2 => n5812, A => n2127, ZN => n3502
                           );
   U1795 : NAND2_X1 port map( A1 => n2111, A2 => n6812, ZN => n2127);
   U1796 : OAI21_X1 port map( B1 => n5504, B2 => n5816, A => n2128, ZN => n3501
                           );
   U1797 : NAND2_X1 port map( A1 => n5812, A2 => n6811, ZN => n2128);
   U1798 : OAI21_X1 port map( B1 => n6073, B2 => n5812, A => n2129, ZN => n3500
                           );
   U1799 : NAND2_X1 port map( A1 => n5812, A2 => n6810, ZN => n2129);
   U1800 : OAI21_X1 port map( B1 => n5498, B2 => n5816, A => n2131, ZN => n3499
                           );
   U1801 : NAND2_X1 port map( A1 => n5812, A2 => n6809, ZN => n2131);
   U1802 : OAI21_X1 port map( B1 => n5495, B2 => n5812, A => n2132, ZN => n3498
                           );
   U1803 : NAND2_X1 port map( A1 => n5812, A2 => n6808, ZN => n2132);
   U1804 : OAI21_X1 port map( B1 => n5492, B2 => n5816, A => n2133, ZN => n3497
                           );
   U1805 : NAND2_X1 port map( A1 => n5812, A2 => n6807, ZN => n2133);
   U1806 : OAI21_X1 port map( B1 => n5489, B2 => n5812, A => n2134, ZN => n3496
                           );
   U1807 : NAND2_X1 port map( A1 => n5812, A2 => n6806, ZN => n2134);
   U1808 : OAI21_X1 port map( B1 => n5486, B2 => n5816, A => n2136, ZN => n3495
                           );
   U1809 : NAND2_X1 port map( A1 => n5812, A2 => n6805, ZN => n2136);
   U1810 : OAI21_X1 port map( B1 => n6067, B2 => n5812, A => n2137, ZN => n3494
                           );
   U1811 : NAND2_X1 port map( A1 => n5812, A2 => n6804, ZN => n2137);
   U1812 : OAI21_X1 port map( B1 => n5480, B2 => n5816, A => n2138, ZN => n3493
                           );
   U1813 : NAND2_X1 port map( A1 => n5816, A2 => n6803, ZN => n2138);
   U1814 : OAI21_X1 port map( B1 => n5477, B2 => n5812, A => n2139, ZN => n3492
                           );
   U1815 : NAND2_X1 port map( A1 => n5816, A2 => n6802, ZN => n2139);
   U1816 : OAI21_X1 port map( B1 => n5474, B2 => n5816, A => n2141, ZN => n3491
                           );
   U1817 : NAND2_X1 port map( A1 => n5816, A2 => n6801, ZN => n2141);
   U1818 : OAI21_X1 port map( B1 => n5471, B2 => n5816, A => n2142, ZN => n3490
                           );
   U1819 : NAND2_X1 port map( A1 => n5816, A2 => n6800, ZN => n2142);
   U1820 : OAI21_X1 port map( B1 => n5468, B2 => n5816, A => n2143, ZN => n3489
                           );
   U1821 : NAND2_X1 port map( A1 => n5812, A2 => n6799, ZN => n2143);
   U1822 : OAI21_X1 port map( B1 => n5465, B2 => n5816, A => n2144, ZN => n3488
                           );
   U1823 : NAND2_X1 port map( A1 => n2111, A2 => n6798, ZN => n2144);
   U1824 : OAI21_X1 port map( B1 => n5462, B2 => n5816, A => n2146, ZN => n3487
                           );
   U1825 : NAND2_X1 port map( A1 => n2111, A2 => n6797, ZN => n2146);
   U1826 : OAI21_X1 port map( B1 => n5459, B2 => n2111, A => n2147, ZN => n3486
                           );
   U1827 : NAND2_X1 port map( A1 => n5816, A2 => n6796, ZN => n2147);
   U1828 : NAND2_X1 port map( A1 => n1556, A2 => n1521, ZN => n2111);
   U1829 : OAI21_X1 port map( B1 => n5552, B2 => n5808, A => n2149, ZN => n3485
                           );
   U1830 : NAND2_X1 port map( A1 => n385, A2 => n2148, ZN => n2149);
   U1831 : OAI21_X1 port map( B1 => n5549, B2 => n5808, A => n2151, ZN => n3484
                           );
   U1832 : NAND2_X1 port map( A1 => n386, A2 => n2148, ZN => n2151);
   U1833 : OAI21_X1 port map( B1 => n5546, B2 => n5808, A => n2152, ZN => n3483
                           );
   U1834 : NAND2_X1 port map( A1 => n387, A2 => n2148, ZN => n2152);
   U1835 : OAI21_X1 port map( B1 => n5543, B2 => n5809, A => n2153, ZN => n3482
                           );
   U1836 : NAND2_X1 port map( A1 => n388, A2 => n2148, ZN => n2153);
   U1837 : OAI21_X1 port map( B1 => n5540, B2 => n5808, A => n2154, ZN => n3481
                           );
   U1838 : NAND2_X1 port map( A1 => n389, A2 => n5809, ZN => n2154);
   U1839 : OAI21_X1 port map( B1 => n5537, B2 => n5808, A => n2156, ZN => n3480
                           );
   U1840 : NAND2_X1 port map( A1 => n390, A2 => n2148, ZN => n2156);
   U1841 : OAI21_X1 port map( B1 => n5534, B2 => n5808, A => n2157, ZN => n3479
                           );
   U1842 : NAND2_X1 port map( A1 => n391, A2 => n2148, ZN => n2157);
   U1843 : OAI21_X1 port map( B1 => n5531, B2 => n5808, A => n2158, ZN => n3478
                           );
   U1844 : NAND2_X1 port map( A1 => n392, A2 => n5808, ZN => n2158);
   U1845 : OAI21_X1 port map( B1 => n5528, B2 => n5808, A => n2159, ZN => n3477
                           );
   U1846 : NAND2_X1 port map( A1 => n393, A2 => n5809, ZN => n2159);
   U1847 : OAI21_X1 port map( B1 => n6081, B2 => n5808, A => n2161, ZN => n3476
                           );
   U1848 : NAND2_X1 port map( A1 => n394, A2 => n5808, ZN => n2161);
   U1849 : OAI21_X1 port map( B1 => n5522, B2 => n5808, A => n2162, ZN => n3475
                           );
   U1850 : NAND2_X1 port map( A1 => n395, A2 => n5809, ZN => n2162);
   U1851 : OAI21_X1 port map( B1 => n5519, B2 => n5808, A => n2163, ZN => n3474
                           );
   U1852 : NAND2_X1 port map( A1 => n396, A2 => n5808, ZN => n2163);
   U1853 : OAI21_X1 port map( B1 => n5516, B2 => n5808, A => n2164, ZN => n3473
                           );
   U1854 : NAND2_X1 port map( A1 => n397, A2 => n5809, ZN => n2164);
   U1855 : OAI21_X1 port map( B1 => n5513, B2 => n5808, A => n2166, ZN => n3472
                           );
   U1856 : NAND2_X1 port map( A1 => n398, A2 => n2148, ZN => n2166);
   U1857 : OAI21_X1 port map( B1 => n5509, B2 => n5808, A => n2167, ZN => n3471
                           );
   U1858 : NAND2_X1 port map( A1 => n399, A2 => n5808, ZN => n2167);
   U1859 : OAI21_X1 port map( B1 => n5506, B2 => n5809, A => n2168, ZN => n3470
                           );
   U1860 : NAND2_X1 port map( A1 => n400, A2 => n5808, ZN => n2168);
   U1861 : OAI21_X1 port map( B1 => n5504, B2 => n5809, A => n2169, ZN => n3469
                           );
   U1862 : NAND2_X1 port map( A1 => n401, A2 => n2148, ZN => n2169);
   U1863 : OAI21_X1 port map( B1 => n6073, B2 => n5809, A => n2171, ZN => n3468
                           );
   U1864 : NAND2_X1 port map( A1 => n402, A2 => n2148, ZN => n2171);
   U1865 : OAI21_X1 port map( B1 => n5498, B2 => n5809, A => n2172, ZN => n3467
                           );
   U1866 : NAND2_X1 port map( A1 => n403, A2 => n2148, ZN => n2172);
   U1867 : OAI21_X1 port map( B1 => n5495, B2 => n5809, A => n2173, ZN => n3466
                           );
   U1868 : NAND2_X1 port map( A1 => n404, A2 => n2148, ZN => n2173);
   U1869 : OAI21_X1 port map( B1 => n5492, B2 => n5809, A => n2174, ZN => n3465
                           );
   U1870 : NAND2_X1 port map( A1 => n405, A2 => n2148, ZN => n2174);
   U1871 : OAI21_X1 port map( B1 => n5489, B2 => n5809, A => n2176, ZN => n3464
                           );
   U1872 : NAND2_X1 port map( A1 => n406, A2 => n2148, ZN => n2176);
   U1873 : OAI21_X1 port map( B1 => n5486, B2 => n5809, A => n2177, ZN => n3463
                           );
   U1874 : NAND2_X1 port map( A1 => n407, A2 => n2148, ZN => n2177);
   U1875 : OAI21_X1 port map( B1 => n6067, B2 => n5809, A => n2178, ZN => n3462
                           );
   U1876 : NAND2_X1 port map( A1 => n408, A2 => n2148, ZN => n2178);
   U1877 : OAI21_X1 port map( B1 => n5480, B2 => n5809, A => n2179, ZN => n3461
                           );
   U1878 : NAND2_X1 port map( A1 => n409, A2 => n2148, ZN => n2179);
   U1879 : OAI21_X1 port map( B1 => n5477, B2 => n5809, A => n2181, ZN => n3460
                           );
   U1880 : NAND2_X1 port map( A1 => n410, A2 => n2148, ZN => n2181);
   U1881 : OAI21_X1 port map( B1 => n5474, B2 => n5809, A => n2182, ZN => n3459
                           );
   U1882 : NAND2_X1 port map( A1 => n411, A2 => n2148, ZN => n2182);
   U1883 : OAI21_X1 port map( B1 => n5471, B2 => n5808, A => n2183, ZN => n3458
                           );
   U1884 : NAND2_X1 port map( A1 => n412, A2 => n2148, ZN => n2183);
   U1885 : OAI21_X1 port map( B1 => n5468, B2 => n5809, A => n2184, ZN => n3457
                           );
   U1886 : NAND2_X1 port map( A1 => n413, A2 => n2148, ZN => n2184);
   U1887 : OAI21_X1 port map( B1 => n5465, B2 => n5808, A => n2186, ZN => n3456
                           );
   U1888 : NAND2_X1 port map( A1 => n414, A2 => n2148, ZN => n2186);
   U1889 : OAI21_X1 port map( B1 => n5462, B2 => n5809, A => n2187, ZN => n3455
                           );
   U1890 : NAND2_X1 port map( A1 => n415, A2 => n2148, ZN => n2187);
   U1891 : OAI21_X1 port map( B1 => n5459, B2 => n5809, A => n2188, ZN => n3454
                           );
   U1892 : NAND2_X1 port map( A1 => n416, A2 => n2148, ZN => n2188);
   U1893 : NAND2_X1 port map( A1 => n1812, A2 => n1556, ZN => n2148);
   U1894 : OAI21_X1 port map( B1 => n5552, B2 => n5804, A => n2191, ZN => n3453
                           );
   U1895 : NAND2_X1 port map( A1 => n417, A2 => n2189, ZN => n2191);
   U1896 : OAI21_X1 port map( B1 => n5549, B2 => n2189, A => n2192, ZN => n3452
                           );
   U1897 : NAND2_X1 port map( A1 => n418, A2 => n2189, ZN => n2192);
   U1898 : OAI21_X1 port map( B1 => n5546, B2 => n5803, A => n2193, ZN => n3451
                           );
   U1899 : NAND2_X1 port map( A1 => n419, A2 => n2189, ZN => n2193);
   U1900 : OAI21_X1 port map( B1 => n5543, B2 => n2189, A => n2194, ZN => n3450
                           );
   U1901 : NAND2_X1 port map( A1 => n420, A2 => n2189, ZN => n2194);
   U1902 : OAI21_X1 port map( B1 => n5540, B2 => n2189, A => n2196, ZN => n3449
                           );
   U1903 : NAND2_X1 port map( A1 => n421, A2 => n5804, ZN => n2196);
   U1904 : OAI21_X1 port map( B1 => n5537, B2 => n5804, A => n2197, ZN => n3448
                           );
   U1905 : NAND2_X1 port map( A1 => n422, A2 => n5804, ZN => n2197);
   U1906 : OAI21_X1 port map( B1 => n5534, B2 => n5803, A => n2198, ZN => n3447
                           );
   U1907 : NAND2_X1 port map( A1 => n423, A2 => n2189, ZN => n2198);
   U1908 : OAI21_X1 port map( B1 => n5531, B2 => n5804, A => n2199, ZN => n3446
                           );
   U1909 : NAND2_X1 port map( A1 => n424, A2 => n2189, ZN => n2199);
   U1910 : OAI21_X1 port map( B1 => n5528, B2 => n5803, A => n2201, ZN => n3445
                           );
   U1911 : NAND2_X1 port map( A1 => n425, A2 => n2189, ZN => n2201);
   U1912 : OAI21_X1 port map( B1 => n6081, B2 => n5804, A => n2202, ZN => n3444
                           );
   U1913 : NAND2_X1 port map( A1 => n426, A2 => n2189, ZN => n2202);
   U1914 : OAI21_X1 port map( B1 => n5522, B2 => n5803, A => n2203, ZN => n3443
                           );
   U1915 : NAND2_X1 port map( A1 => n427, A2 => n2189, ZN => n2203);
   U1916 : OAI21_X1 port map( B1 => n5519, B2 => n5804, A => n2204, ZN => n3442
                           );
   U1917 : NAND2_X1 port map( A1 => n428, A2 => n2189, ZN => n2204);
   U1918 : OAI21_X1 port map( B1 => n5516, B2 => n5803, A => n2206, ZN => n3441
                           );
   U1919 : NAND2_X1 port map( A1 => n429, A2 => n2189, ZN => n2206);
   U1920 : OAI21_X1 port map( B1 => n5513, B2 => n5804, A => n2207, ZN => n3440
                           );
   U1921 : NAND2_X1 port map( A1 => n430, A2 => n2189, ZN => n2207);
   U1922 : OAI21_X1 port map( B1 => n5509, B2 => n2189, A => n2208, ZN => n3439
                           );
   U1923 : NAND2_X1 port map( A1 => n431, A2 => n2189, ZN => n2208);
   U1924 : OAI21_X1 port map( B1 => n6075, B2 => n5803, A => n2209, ZN => n3438
                           );
   U1925 : NAND2_X1 port map( A1 => n432, A2 => n5804, ZN => n2209);
   U1926 : OAI21_X1 port map( B1 => n6074, B2 => n5803, A => n2211, ZN => n3437
                           );
   U1927 : NAND2_X1 port map( A1 => n433, A2 => n5803, ZN => n2211);
   U1928 : OAI21_X1 port map( B1 => n5499, B2 => n5803, A => n2212, ZN => n3436
                           );
   U1929 : NAND2_X1 port map( A1 => n434, A2 => n5804, ZN => n2212);
   U1930 : OAI21_X1 port map( B1 => n6072, B2 => n5803, A => n2213, ZN => n3435
                           );
   U1931 : NAND2_X1 port map( A1 => n435, A2 => n5804, ZN => n2213);
   U1932 : OAI21_X1 port map( B1 => n6071, B2 => n5803, A => n2214, ZN => n3434
                           );
   U1933 : NAND2_X1 port map( A1 => n436, A2 => n5804, ZN => n2214);
   U1934 : OAI21_X1 port map( B1 => n6070, B2 => n5803, A => n2216, ZN => n3433
                           );
   U1935 : NAND2_X1 port map( A1 => n437, A2 => n5804, ZN => n2216);
   U1936 : OAI21_X1 port map( B1 => n6069, B2 => n5803, A => n2217, ZN => n3432
                           );
   U1937 : NAND2_X1 port map( A1 => n438, A2 => n5804, ZN => n2217);
   U1938 : OAI21_X1 port map( B1 => n6068, B2 => n5803, A => n2218, ZN => n3431
                           );
   U1939 : NAND2_X1 port map( A1 => n439, A2 => n5804, ZN => n2218);
   U1940 : OAI21_X1 port map( B1 => n5481, B2 => n5803, A => n2219, ZN => n3430
                           );
   U1941 : NAND2_X1 port map( A1 => n440, A2 => n5804, ZN => n2219);
   U1942 : OAI21_X1 port map( B1 => n6066, B2 => n5803, A => n2221, ZN => n3429
                           );
   U1943 : NAND2_X1 port map( A1 => n441, A2 => n2189, ZN => n2221);
   U1944 : OAI21_X1 port map( B1 => n6065, B2 => n5803, A => n2222, ZN => n3428
                           );
   U1945 : NAND2_X1 port map( A1 => n442, A2 => n2189, ZN => n2222);
   U1946 : OAI21_X1 port map( B1 => n6064, B2 => n5803, A => n2223, ZN => n3427
                           );
   U1947 : NAND2_X1 port map( A1 => n443, A2 => n2189, ZN => n2223);
   U1948 : OAI21_X1 port map( B1 => n6063, B2 => n5804, A => n2224, ZN => n3426
                           );
   U1949 : NAND2_X1 port map( A1 => n444, A2 => n2189, ZN => n2224);
   U1950 : OAI21_X1 port map( B1 => n6062, B2 => n5804, A => n2226, ZN => n3425
                           );
   U1951 : NAND2_X1 port map( A1 => n445, A2 => n2189, ZN => n2226);
   U1952 : OAI21_X1 port map( B1 => n6061, B2 => n5804, A => n2227, ZN => n3424
                           );
   U1953 : NAND2_X1 port map( A1 => n446, A2 => n2189, ZN => n2227);
   U1954 : OAI21_X1 port map( B1 => n6060, B2 => n5804, A => n2228, ZN => n3423
                           );
   U1955 : NAND2_X1 port map( A1 => n447, A2 => n5803, ZN => n2228);
   U1956 : OAI21_X1 port map( B1 => n6059, B2 => n2189, A => n2229, ZN => n3422
                           );
   U1957 : NAND2_X1 port map( A1 => n448, A2 => n5803, ZN => n2229);
   U1958 : NAND2_X1 port map( A1 => n1778, A2 => n1556, ZN => n2189);
   U1959 : OAI21_X1 port map( B1 => n6090, B2 => n5793, A => n2232, ZN => n3421
                           );
   U1960 : NAND2_X1 port map( A1 => n545, A2 => n5793, ZN => n2232);
   U1961 : OAI21_X1 port map( B1 => n6089, B2 => n5795, A => n2233, ZN => n3420
                           );
   U1962 : NAND2_X1 port map( A1 => n546, A2 => n5793, ZN => n2233);
   U1963 : OAI21_X1 port map( B1 => n6088, B2 => n2231, A => n2234, ZN => n3419
                           );
   U1964 : NAND2_X1 port map( A1 => n547, A2 => n5793, ZN => n2234);
   U1965 : OAI21_X1 port map( B1 => n6087, B2 => n5795, A => n2236, ZN => n3418
                           );
   U1966 : NAND2_X1 port map( A1 => n548, A2 => n5793, ZN => n2236);
   U1967 : OAI21_X1 port map( B1 => n6086, B2 => n5795, A => n2237, ZN => n3417
                           );
   U1968 : NAND2_X1 port map( A1 => n549, A2 => n5795, ZN => n2237);
   U1969 : OAI21_X1 port map( B1 => n6085, B2 => n2231, A => n2238, ZN => n3416
                           );
   U1970 : NAND2_X1 port map( A1 => n550, A2 => n5795, ZN => n2238);
   U1971 : OAI21_X1 port map( B1 => n6084, B2 => n2231, A => n2239, ZN => n3415
                           );
   U1972 : NAND2_X1 port map( A1 => n551, A2 => n5793, ZN => n2239);
   U1973 : OAI21_X1 port map( B1 => n6083, B2 => n2231, A => n2241, ZN => n3414
                           );
   U1974 : NAND2_X1 port map( A1 => n552, A2 => n5795, ZN => n2241);
   U1975 : OAI21_X1 port map( B1 => n6082, B2 => n2231, A => n2242, ZN => n3413
                           );
   U1976 : NAND2_X1 port map( A1 => n553, A2 => n5795, ZN => n2242);
   U1977 : OAI21_X1 port map( B1 => n5523, B2 => n2231, A => n2243, ZN => n3412
                           );
   U1978 : NAND2_X1 port map( A1 => n554, A2 => n5795, ZN => n2243);
   U1979 : OAI21_X1 port map( B1 => n6080, B2 => n2231, A => n2244, ZN => n3411
                           );
   U1980 : NAND2_X1 port map( A1 => n555, A2 => n5795, ZN => n2244);
   U1981 : OAI21_X1 port map( B1 => n6079, B2 => n2231, A => n2246, ZN => n3410
                           );
   U1982 : NAND2_X1 port map( A1 => n556, A2 => n5795, ZN => n2246);
   U1983 : OAI21_X1 port map( B1 => n6078, B2 => n2231, A => n2247, ZN => n3409
                           );
   U1984 : NAND2_X1 port map( A1 => n557, A2 => n5795, ZN => n2247);
   U1985 : OAI21_X1 port map( B1 => n6077, B2 => n2231, A => n2248, ZN => n3408
                           );
   U1986 : NAND2_X1 port map( A1 => n558, A2 => n5795, ZN => n2248);
   U1987 : OAI21_X1 port map( B1 => n6076, B2 => n2231, A => n2249, ZN => n3407
                           );
   U1988 : NAND2_X1 port map( A1 => n559, A2 => n5795, ZN => n2249);
   U1989 : OAI21_X1 port map( B1 => n6075, B2 => n2231, A => n2251, ZN => n3406
                           );
   U1990 : NAND2_X1 port map( A1 => n560, A2 => n5795, ZN => n2251);
   U1991 : OAI21_X1 port map( B1 => n6074, B2 => n2231, A => n2252, ZN => n3405
                           );
   U1992 : NAND2_X1 port map( A1 => n561, A2 => n5793, ZN => n2252);
   U1993 : OAI21_X1 port map( B1 => n5499, B2 => n2231, A => n2253, ZN => n3404
                           );
   U1994 : NAND2_X1 port map( A1 => n562, A2 => n5795, ZN => n2253);
   U1995 : OAI21_X1 port map( B1 => n6072, B2 => n2231, A => n2254, ZN => n3403
                           );
   U1996 : NAND2_X1 port map( A1 => n563, A2 => n5793, ZN => n2254);
   U1997 : OAI21_X1 port map( B1 => n6071, B2 => n2231, A => n2256, ZN => n3402
                           );
   U1998 : NAND2_X1 port map( A1 => n564, A2 => n5795, ZN => n2256);
   U1999 : OAI21_X1 port map( B1 => n6070, B2 => n2231, A => n2257, ZN => n3401
                           );
   U2000 : NAND2_X1 port map( A1 => n565, A2 => n5793, ZN => n2257);
   U2001 : OAI21_X1 port map( B1 => n6069, B2 => n2231, A => n2258, ZN => n3400
                           );
   U2002 : NAND2_X1 port map( A1 => n566, A2 => n5795, ZN => n2258);
   U2003 : OAI21_X1 port map( B1 => n6068, B2 => n2231, A => n2259, ZN => n3399
                           );
   U2004 : NAND2_X1 port map( A1 => n567, A2 => n5793, ZN => n2259);
   U2005 : OAI21_X1 port map( B1 => n5481, B2 => n2231, A => n2261, ZN => n3398
                           );
   U2006 : NAND2_X1 port map( A1 => n568, A2 => n5795, ZN => n2261);
   U2007 : OAI21_X1 port map( B1 => n6066, B2 => n5795, A => n2262, ZN => n3397
                           );
   U2008 : NAND2_X1 port map( A1 => n569, A2 => n5793, ZN => n2262);
   U2009 : OAI21_X1 port map( B1 => n6065, B2 => n2231, A => n2263, ZN => n3396
                           );
   U2010 : NAND2_X1 port map( A1 => n570, A2 => n5793, ZN => n2263);
   U2011 : OAI21_X1 port map( B1 => n6064, B2 => n2231, A => n2264, ZN => n3395
                           );
   U2012 : NAND2_X1 port map( A1 => n571, A2 => n5793, ZN => n2264);
   U2013 : OAI21_X1 port map( B1 => n6063, B2 => n2231, A => n2266, ZN => n3394
                           );
   U2014 : NAND2_X1 port map( A1 => n572, A2 => n5793, ZN => n2266);
   U2015 : OAI21_X1 port map( B1 => n6062, B2 => n2231, A => n2267, ZN => n3393
                           );
   U2016 : NAND2_X1 port map( A1 => n573, A2 => n5793, ZN => n2267);
   U2017 : OAI21_X1 port map( B1 => n6061, B2 => n5793, A => n2268, ZN => n3392
                           );
   U2018 : NAND2_X1 port map( A1 => n574, A2 => n5793, ZN => n2268);
   U2019 : OAI21_X1 port map( B1 => n6060, B2 => n5793, A => n2269, ZN => n3391
                           );
   U2020 : NAND2_X1 port map( A1 => n575, A2 => n5793, ZN => n2269);
   U2021 : OAI21_X1 port map( B1 => n6059, B2 => n5795, A => n2271, ZN => n3390
                           );
   U2022 : NAND2_X1 port map( A1 => n576, A2 => n5793, ZN => n2271);
   U2023 : NAND2_X1 port map( A1 => n2110, A2 => n1556, ZN => n2231);
   U2024 : NOR2_X1 port map( A1 => n2272, A2 => n6048, ZN => n1556);
   U2025 : OR2_X1 port map( A1 => ADD_WR(4), A2 => n2273, ZN => n2272);
   U2026 : OAI21_X1 port map( B1 => n6090, B2 => n5790, A => n2275, ZN => n3389
                           );
   U2027 : NAND2_X1 port map( A1 => n449, A2 => n2274, ZN => n2275);
   U2028 : OAI21_X1 port map( B1 => n6089, B2 => n5790, A => n2276, ZN => n3388
                           );
   U2029 : NAND2_X1 port map( A1 => n450, A2 => n2274, ZN => n2276);
   U2030 : OAI21_X1 port map( B1 => n6088, B2 => n5790, A => n2277, ZN => n3387
                           );
   U2031 : NAND2_X1 port map( A1 => n451, A2 => n2274, ZN => n2277);
   U2032 : OAI21_X1 port map( B1 => n6087, B2 => n5791, A => n2278, ZN => n3386
                           );
   U2033 : NAND2_X1 port map( A1 => n452, A2 => n2274, ZN => n2278);
   U2034 : OAI21_X1 port map( B1 => n6086, B2 => n5790, A => n2279, ZN => n3385
                           );
   U2035 : NAND2_X1 port map( A1 => n453, A2 => n5791, ZN => n2279);
   U2036 : OAI21_X1 port map( B1 => n6085, B2 => n5790, A => n2280, ZN => n3384
                           );
   U2037 : NAND2_X1 port map( A1 => n454, A2 => n2274, ZN => n2280);
   U2038 : OAI21_X1 port map( B1 => n6084, B2 => n5790, A => n2281, ZN => n3383
                           );
   U2039 : NAND2_X1 port map( A1 => n455, A2 => n2274, ZN => n2281);
   U2040 : OAI21_X1 port map( B1 => n6083, B2 => n5790, A => n2282, ZN => n3382
                           );
   U2041 : NAND2_X1 port map( A1 => n456, A2 => n5790, ZN => n2282);
   U2042 : OAI21_X1 port map( B1 => n6082, B2 => n5790, A => n2283, ZN => n3381
                           );
   U2043 : NAND2_X1 port map( A1 => n457, A2 => n5791, ZN => n2283);
   U2044 : OAI21_X1 port map( B1 => n5523, B2 => n5790, A => n2284, ZN => n3380
                           );
   U2045 : NAND2_X1 port map( A1 => n458, A2 => n5790, ZN => n2284);
   U2046 : OAI21_X1 port map( B1 => n6080, B2 => n5790, A => n2285, ZN => n3379
                           );
   U2047 : NAND2_X1 port map( A1 => n459, A2 => n5791, ZN => n2285);
   U2048 : OAI21_X1 port map( B1 => n6079, B2 => n5790, A => n2286, ZN => n3378
                           );
   U2049 : NAND2_X1 port map( A1 => n460, A2 => n5790, ZN => n2286);
   U2050 : OAI21_X1 port map( B1 => n6078, B2 => n5790, A => n2287, ZN => n3377
                           );
   U2051 : NAND2_X1 port map( A1 => n461, A2 => n5791, ZN => n2287);
   U2052 : OAI21_X1 port map( B1 => n6077, B2 => n5790, A => n2288, ZN => n3376
                           );
   U2053 : NAND2_X1 port map( A1 => n462, A2 => n2274, ZN => n2288);
   U2054 : OAI21_X1 port map( B1 => n6076, B2 => n5790, A => n2289, ZN => n3375
                           );
   U2055 : NAND2_X1 port map( A1 => n463, A2 => n5790, ZN => n2289);
   U2056 : OAI21_X1 port map( B1 => n6075, B2 => n5791, A => n2290, ZN => n3374
                           );
   U2057 : NAND2_X1 port map( A1 => n464, A2 => n5790, ZN => n2290);
   U2058 : OAI21_X1 port map( B1 => n6074, B2 => n5791, A => n2291, ZN => n3373
                           );
   U2059 : NAND2_X1 port map( A1 => n465, A2 => n2274, ZN => n2291);
   U2060 : OAI21_X1 port map( B1 => n5499, B2 => n5791, A => n2292, ZN => n3372
                           );
   U2061 : NAND2_X1 port map( A1 => n466, A2 => n2274, ZN => n2292);
   U2062 : OAI21_X1 port map( B1 => n6072, B2 => n5791, A => n2293, ZN => n3371
                           );
   U2063 : NAND2_X1 port map( A1 => n467, A2 => n2274, ZN => n2293);
   U2064 : OAI21_X1 port map( B1 => n6071, B2 => n5791, A => n2294, ZN => n3370
                           );
   U2065 : NAND2_X1 port map( A1 => n468, A2 => n2274, ZN => n2294);
   U2066 : OAI21_X1 port map( B1 => n6070, B2 => n5791, A => n2295, ZN => n3369
                           );
   U2067 : NAND2_X1 port map( A1 => n469, A2 => n2274, ZN => n2295);
   U2068 : OAI21_X1 port map( B1 => n6069, B2 => n5791, A => n2296, ZN => n3368
                           );
   U2069 : NAND2_X1 port map( A1 => n470, A2 => n2274, ZN => n2296);
   U2070 : OAI21_X1 port map( B1 => n6068, B2 => n5791, A => n2297, ZN => n3367
                           );
   U2071 : NAND2_X1 port map( A1 => n471, A2 => n2274, ZN => n2297);
   U2072 : OAI21_X1 port map( B1 => n5481, B2 => n5791, A => n2298, ZN => n3366
                           );
   U2073 : NAND2_X1 port map( A1 => n472, A2 => n2274, ZN => n2298);
   U2074 : OAI21_X1 port map( B1 => n6066, B2 => n5791, A => n2299, ZN => n3365
                           );
   U2075 : NAND2_X1 port map( A1 => n473, A2 => n2274, ZN => n2299);
   U2076 : OAI21_X1 port map( B1 => n6065, B2 => n5791, A => n2300, ZN => n3364
                           );
   U2077 : NAND2_X1 port map( A1 => n474, A2 => n2274, ZN => n2300);
   U2078 : OAI21_X1 port map( B1 => n6064, B2 => n5791, A => n2301, ZN => n3363
                           );
   U2079 : NAND2_X1 port map( A1 => n475, A2 => n2274, ZN => n2301);
   U2080 : OAI21_X1 port map( B1 => n6063, B2 => n5790, A => n2302, ZN => n3362
                           );
   U2081 : NAND2_X1 port map( A1 => n476, A2 => n2274, ZN => n2302);
   U2082 : OAI21_X1 port map( B1 => n6062, B2 => n5791, A => n2303, ZN => n3361
                           );
   U2083 : NAND2_X1 port map( A1 => n477, A2 => n2274, ZN => n2303);
   U2084 : OAI21_X1 port map( B1 => n6061, B2 => n5790, A => n2304, ZN => n3360
                           );
   U2085 : NAND2_X1 port map( A1 => n478, A2 => n2274, ZN => n2304);
   U2086 : OAI21_X1 port map( B1 => n6060, B2 => n5791, A => n2305, ZN => n3359
                           );
   U2087 : NAND2_X1 port map( A1 => n479, A2 => n2274, ZN => n2305);
   U2088 : OAI21_X1 port map( B1 => n6059, B2 => n5791, A => n2306, ZN => n3358
                           );
   U2089 : NAND2_X1 port map( A1 => n480, A2 => n2274, ZN => n2306);
   U2090 : NAND2_X1 port map( A1 => n1658, A2 => n1520, ZN => n2274);
   U2092 : NOR2_X1 port map( A1 => n6050, A2 => n6049, ZN => n2307);
   U2093 : OAI21_X1 port map( B1 => n6090, B2 => n5785, A => n2309, ZN => n3357
                           );
   U2094 : NAND2_X1 port map( A1 => n2308, A2 => n6795, ZN => n2309);
   U2095 : OAI21_X1 port map( B1 => n6089, B2 => n2308, A => n2310, ZN => n3356
                           );
   U2096 : NAND2_X1 port map( A1 => n2308, A2 => n6794, ZN => n2310);
   U2097 : OAI21_X1 port map( B1 => n6088, B2 => n5786, A => n2311, ZN => n3355
                           );
   U2098 : NAND2_X1 port map( A1 => n2308, A2 => n6793, ZN => n2311);
   U2099 : OAI21_X1 port map( B1 => n6087, B2 => n2308, A => n2312, ZN => n3354
                           );
   U2100 : NAND2_X1 port map( A1 => n2308, A2 => n6792, ZN => n2312);
   U2101 : OAI21_X1 port map( B1 => n6086, B2 => n2308, A => n2313, ZN => n3353
                           );
   U2102 : NAND2_X1 port map( A1 => n5786, A2 => n6791, ZN => n2313);
   U2103 : OAI21_X1 port map( B1 => n6085, B2 => n5785, A => n2314, ZN => n3352
                           );
   U2104 : NAND2_X1 port map( A1 => n5786, A2 => n6790, ZN => n2314);
   U2105 : OAI21_X1 port map( B1 => n6084, B2 => n5786, A => n2315, ZN => n3351
                           );
   U2106 : NAND2_X1 port map( A1 => n2308, A2 => n6789, ZN => n2315);
   U2107 : OAI21_X1 port map( B1 => n6083, B2 => n5785, A => n2316, ZN => n3350
                           );
   U2108 : NAND2_X1 port map( A1 => n2308, A2 => n6788, ZN => n2316);
   U2109 : OAI21_X1 port map( B1 => n6082, B2 => n5786, A => n2317, ZN => n3349
                           );
   U2110 : NAND2_X1 port map( A1 => n2308, A2 => n6787, ZN => n2317);
   U2111 : OAI21_X1 port map( B1 => n5523, B2 => n5785, A => n2318, ZN => n3348
                           );
   U2112 : NAND2_X1 port map( A1 => n2308, A2 => n6786, ZN => n2318);
   U2113 : OAI21_X1 port map( B1 => n6080, B2 => n5786, A => n2319, ZN => n3347
                           );
   U2114 : NAND2_X1 port map( A1 => n2308, A2 => n6785, ZN => n2319);
   U2115 : OAI21_X1 port map( B1 => n6079, B2 => n5785, A => n2320, ZN => n3346
                           );
   U2116 : NAND2_X1 port map( A1 => n2308, A2 => n6784, ZN => n2320);
   U2117 : OAI21_X1 port map( B1 => n6078, B2 => n5786, A => n2321, ZN => n3345
                           );
   U2118 : NAND2_X1 port map( A1 => n2308, A2 => n6783, ZN => n2321);
   U2119 : OAI21_X1 port map( B1 => n6077, B2 => n2308, A => n2322, ZN => n3344
                           );
   U2120 : NAND2_X1 port map( A1 => n5786, A2 => n6782, ZN => n2322);
   U2121 : OAI21_X1 port map( B1 => n6076, B2 => n2308, A => n2323, ZN => n3343
                           );
   U2122 : NAND2_X1 port map( A1 => n2308, A2 => n6781, ZN => n2323);
   U2123 : OAI21_X1 port map( B1 => n6075, B2 => n5785, A => n2324, ZN => n3342
                           );
   U2124 : NAND2_X1 port map( A1 => n5785, A2 => n6780, ZN => n2324);
   U2125 : OAI21_X1 port map( B1 => n6074, B2 => n5785, A => n2325, ZN => n3341
                           );
   U2126 : NAND2_X1 port map( A1 => n5785, A2 => n6779, ZN => n2325);
   U2127 : OAI21_X1 port map( B1 => n5499, B2 => n5785, A => n2326, ZN => n3340
                           );
   U2128 : NAND2_X1 port map( A1 => n5786, A2 => n6778, ZN => n2326);
   U2129 : OAI21_X1 port map( B1 => n6072, B2 => n5785, A => n2327, ZN => n3339
                           );
   U2130 : NAND2_X1 port map( A1 => n5786, A2 => n6777, ZN => n2327);
   U2131 : OAI21_X1 port map( B1 => n6071, B2 => n5785, A => n2328, ZN => n3338
                           );
   U2132 : NAND2_X1 port map( A1 => n5786, A2 => n6776, ZN => n2328);
   U2133 : OAI21_X1 port map( B1 => n6070, B2 => n5785, A => n2329, ZN => n3337
                           );
   U2134 : NAND2_X1 port map( A1 => n5786, A2 => n6775, ZN => n2329);
   U2135 : OAI21_X1 port map( B1 => n6069, B2 => n5785, A => n2330, ZN => n3336
                           );
   U2136 : NAND2_X1 port map( A1 => n5786, A2 => n6774, ZN => n2330);
   U2137 : OAI21_X1 port map( B1 => n6068, B2 => n5785, A => n2331, ZN => n3335
                           );
   U2138 : NAND2_X1 port map( A1 => n5786, A2 => n6773, ZN => n2331);
   U2139 : OAI21_X1 port map( B1 => n5481, B2 => n5785, A => n2332, ZN => n3334
                           );
   U2140 : NAND2_X1 port map( A1 => n5786, A2 => n6772, ZN => n2332);
   U2141 : OAI21_X1 port map( B1 => n6066, B2 => n5785, A => n2333, ZN => n3333
                           );
   U2142 : NAND2_X1 port map( A1 => n2308, A2 => n6771, ZN => n2333);
   U2143 : OAI21_X1 port map( B1 => n6065, B2 => n5785, A => n2334, ZN => n3332
                           );
   U2144 : NAND2_X1 port map( A1 => n2308, A2 => n6770, ZN => n2334);
   U2145 : OAI21_X1 port map( B1 => n6064, B2 => n5785, A => n2335, ZN => n3331
                           );
   U2146 : NAND2_X1 port map( A1 => n2308, A2 => n6769, ZN => n2335);
   U2147 : OAI21_X1 port map( B1 => n6063, B2 => n5786, A => n2336, ZN => n3330
                           );
   U2148 : NAND2_X1 port map( A1 => n2308, A2 => n6768, ZN => n2336);
   U2149 : OAI21_X1 port map( B1 => n6062, B2 => n5786, A => n2337, ZN => n3329
                           );
   U2150 : NAND2_X1 port map( A1 => n5786, A2 => n6767, ZN => n2337);
   U2151 : OAI21_X1 port map( B1 => n6061, B2 => n5786, A => n2338, ZN => n3328
                           );
   U2152 : NAND2_X1 port map( A1 => n2308, A2 => n6766, ZN => n2338);
   U2153 : OAI21_X1 port map( B1 => n6060, B2 => n5786, A => n2339, ZN => n3327
                           );
   U2154 : NAND2_X1 port map( A1 => n2308, A2 => n6765, ZN => n2339);
   U2155 : OAI21_X1 port map( B1 => n6059, B2 => n2308, A => n2340, ZN => n3326
                           );
   U2156 : NAND2_X1 port map( A1 => n5785, A2 => n6764, ZN => n2340);
   U2157 : NAND2_X1 port map( A1 => n1624, A2 => n1520, ZN => n2308);
   U2159 : NOR2_X1 port map( A1 => ADD_WR(0), A2 => n6049, ZN => n2341);
   U2160 : OAI21_X1 port map( B1 => n6090, B2 => n2342, A => n2343, ZN => n3325
                           );
   U2161 : NAND2_X1 port map( A1 => n577, A2 => n5775, ZN => n2343);
   U2162 : OAI21_X1 port map( B1 => n6089, B2 => n5777, A => n2344, ZN => n3324
                           );
   U2163 : NAND2_X1 port map( A1 => n578, A2 => n5775, ZN => n2344);
   U2164 : OAI21_X1 port map( B1 => n6088, B2 => n2342, A => n2345, ZN => n3323
                           );
   U2165 : NAND2_X1 port map( A1 => n579, A2 => n5775, ZN => n2345);
   U2166 : OAI21_X1 port map( B1 => n6087, B2 => n5777, A => n2346, ZN => n3322
                           );
   U2167 : NAND2_X1 port map( A1 => n580, A2 => n5775, ZN => n2346);
   U2168 : OAI21_X1 port map( B1 => n6086, B2 => n5777, A => n2347, ZN => n3321
                           );
   U2169 : NAND2_X1 port map( A1 => n581, A2 => n5775, ZN => n2347);
   U2170 : OAI21_X1 port map( B1 => n6085, B2 => n2342, A => n2348, ZN => n3320
                           );
   U2171 : NAND2_X1 port map( A1 => n582, A2 => n5775, ZN => n2348);
   U2172 : OAI21_X1 port map( B1 => n6084, B2 => n2342, A => n2349, ZN => n3319
                           );
   U2173 : NAND2_X1 port map( A1 => n583, A2 => n5777, ZN => n2349);
   U2174 : OAI21_X1 port map( B1 => n6083, B2 => n2342, A => n2350, ZN => n3318
                           );
   U2175 : NAND2_X1 port map( A1 => n584, A2 => n5777, ZN => n2350);
   U2176 : OAI21_X1 port map( B1 => n6082, B2 => n2342, A => n2351, ZN => n3317
                           );
   U2177 : NAND2_X1 port map( A1 => n585, A2 => n5777, ZN => n2351);
   U2178 : OAI21_X1 port map( B1 => n5523, B2 => n2342, A => n2353, ZN => n3316
                           );
   U2179 : NAND2_X1 port map( A1 => n586, A2 => n5777, ZN => n2353);
   U2180 : OAI21_X1 port map( B1 => n6080, B2 => n2342, A => n2354, ZN => n3315
                           );
   U2181 : NAND2_X1 port map( A1 => n587, A2 => n5777, ZN => n2354);
   U2182 : OAI21_X1 port map( B1 => n6079, B2 => n2342, A => n2356, ZN => n3314
                           );
   U2183 : NAND2_X1 port map( A1 => n588, A2 => n5777, ZN => n2356);
   U2184 : OAI21_X1 port map( B1 => n6078, B2 => n2342, A => n2357, ZN => n3313
                           );
   U2185 : NAND2_X1 port map( A1 => n589, A2 => n5777, ZN => n2357);
   U2186 : OAI21_X1 port map( B1 => n6077, B2 => n2342, A => n2359, ZN => n3312
                           );
   U2187 : NAND2_X1 port map( A1 => n590, A2 => n5775, ZN => n2359);
   U2188 : OAI21_X1 port map( B1 => n6076, B2 => n2342, A => n2360, ZN => n3311
                           );
   U2189 : NAND2_X1 port map( A1 => n591, A2 => n5777, ZN => n2360);
   U2190 : OAI21_X1 port map( B1 => n6075, B2 => n2342, A => n2362, ZN => n3310
                           );
   U2191 : NAND2_X1 port map( A1 => n592, A2 => n5777, ZN => n2362);
   U2192 : OAI21_X1 port map( B1 => n6074, B2 => n2342, A => n2363, ZN => n3309
                           );
   U2193 : NAND2_X1 port map( A1 => n593, A2 => n5777, ZN => n2363);
   U2194 : OAI21_X1 port map( B1 => n5499, B2 => n2342, A => n2365, ZN => n3308
                           );
   U2195 : NAND2_X1 port map( A1 => n594, A2 => n5775, ZN => n2365);
   U2196 : OAI21_X1 port map( B1 => n6072, B2 => n2342, A => n2366, ZN => n3307
                           );
   U2197 : NAND2_X1 port map( A1 => n595, A2 => n5777, ZN => n2366);
   U2198 : OAI21_X1 port map( B1 => n6071, B2 => n2342, A => n2368, ZN => n3306
                           );
   U2199 : NAND2_X1 port map( A1 => n596, A2 => n5775, ZN => n2368);
   U2200 : OAI21_X1 port map( B1 => n6070, B2 => n2342, A => n2369, ZN => n3305
                           );
   U2201 : NAND2_X1 port map( A1 => n597, A2 => n5777, ZN => n2369);
   U2202 : OAI21_X1 port map( B1 => n6069, B2 => n2342, A => n2371, ZN => n3304
                           );
   U2203 : NAND2_X1 port map( A1 => n598, A2 => n5775, ZN => n2371);
   U2204 : OAI21_X1 port map( B1 => n6068, B2 => n5777, A => n2372, ZN => n3303
                           );
   U2205 : NAND2_X1 port map( A1 => n599, A2 => n5777, ZN => n2372);
   U2206 : OAI21_X1 port map( B1 => n5481, B2 => n5775, A => n2374, ZN => n3302
                           );
   U2207 : NAND2_X1 port map( A1 => n600, A2 => n5775, ZN => n2374);
   U2208 : OAI21_X1 port map( B1 => n6066, B2 => n5777, A => n2375, ZN => n3301
                           );
   U2209 : NAND2_X1 port map( A1 => n601, A2 => n5775, ZN => n2375);
   U2210 : OAI21_X1 port map( B1 => n6065, B2 => n2342, A => n2377, ZN => n3300
                           );
   U2211 : NAND2_X1 port map( A1 => n602, A2 => n5775, ZN => n2377);
   U2212 : OAI21_X1 port map( B1 => n6064, B2 => n2342, A => n2378, ZN => n3299
                           );
   U2213 : NAND2_X1 port map( A1 => n603, A2 => n5775, ZN => n2378);
   U2214 : OAI21_X1 port map( B1 => n6063, B2 => n2342, A => n2380, ZN => n3298
                           );
   U2215 : NAND2_X1 port map( A1 => n604, A2 => n5775, ZN => n2380);
   U2216 : OAI21_X1 port map( B1 => n6062, B2 => n2342, A => n2381, ZN => n3297
                           );
   U2217 : NAND2_X1 port map( A1 => n605, A2 => n5775, ZN => n2381);
   U2218 : OAI21_X1 port map( B1 => n6061, B2 => n2342, A => n2383, ZN => n3296
                           );
   U2219 : NAND2_X1 port map( A1 => n606, A2 => n5775, ZN => n2383);
   U2220 : OAI21_X1 port map( B1 => n6060, B2 => n5777, A => n2384, ZN => n3295
                           );
   U2221 : NAND2_X1 port map( A1 => n607, A2 => n5775, ZN => n2384);
   U2222 : OAI21_X1 port map( B1 => n6059, B2 => n5777, A => n2385, ZN => n3294
                           );
   U2223 : NAND2_X1 port map( A1 => n608, A2 => n5775, ZN => n2385);
   U2224 : NAND2_X1 port map( A1 => n1590, A2 => n1520, ZN => n2342);
   U2225 : OAI21_X1 port map( B1 => n6090, B2 => n5773, A => n2387, ZN => n3293
                           );
   U2226 : NAND2_X1 port map( A1 => n2386, A2 => n6970, ZN => n2387);
   U2227 : OAI21_X1 port map( B1 => n6089, B2 => n2386, A => n2388, ZN => n3292
                           );
   U2228 : NAND2_X1 port map( A1 => n2386, A2 => n6969, ZN => n2388);
   U2229 : OAI21_X1 port map( B1 => n6088, B2 => n5774, A => n2389, ZN => n3291
                           );
   U2230 : NAND2_X1 port map( A1 => n2386, A2 => n6968, ZN => n2389);
   U2231 : OAI21_X1 port map( B1 => n6087, B2 => n2386, A => n2390, ZN => n3290
                           );
   U2232 : NAND2_X1 port map( A1 => n2386, A2 => n6967, ZN => n2390);
   U2233 : OAI21_X1 port map( B1 => n6086, B2 => n2386, A => n2391, ZN => n3289
                           );
   U2234 : NAND2_X1 port map( A1 => n5774, A2 => n6966, ZN => n2391);
   U2235 : OAI21_X1 port map( B1 => n6085, B2 => n5773, A => n2392, ZN => n3288
                           );
   U2236 : NAND2_X1 port map( A1 => n5774, A2 => n6965, ZN => n2392);
   U2237 : OAI21_X1 port map( B1 => n6084, B2 => n5774, A => n2393, ZN => n3287
                           );
   U2238 : NAND2_X1 port map( A1 => n2386, A2 => n6964, ZN => n2393);
   U2239 : OAI21_X1 port map( B1 => n6083, B2 => n5773, A => n2394, ZN => n3286
                           );
   U2240 : NAND2_X1 port map( A1 => n2386, A2 => n6963, ZN => n2394);
   U2241 : OAI21_X1 port map( B1 => n6082, B2 => n5774, A => n2395, ZN => n3285
                           );
   U2242 : NAND2_X1 port map( A1 => n2386, A2 => n6962, ZN => n2395);
   U2243 : OAI21_X1 port map( B1 => n5523, B2 => n5773, A => n2396, ZN => n3284
                           );
   U2244 : NAND2_X1 port map( A1 => n2386, A2 => n6961, ZN => n2396);
   U2245 : OAI21_X1 port map( B1 => n6080, B2 => n5774, A => n2397, ZN => n3283
                           );
   U2246 : NAND2_X1 port map( A1 => n2386, A2 => n6960, ZN => n2397);
   U2247 : OAI21_X1 port map( B1 => n6079, B2 => n5773, A => n2398, ZN => n3282
                           );
   U2248 : NAND2_X1 port map( A1 => n2386, A2 => n6959, ZN => n2398);
   U2249 : OAI21_X1 port map( B1 => n6078, B2 => n5774, A => n2399, ZN => n3281
                           );
   U2250 : NAND2_X1 port map( A1 => n2386, A2 => n6958, ZN => n2399);
   U2251 : OAI21_X1 port map( B1 => n6077, B2 => n2386, A => n2400, ZN => n3280
                           );
   U2252 : NAND2_X1 port map( A1 => n5774, A2 => n6957, ZN => n2400);
   U2253 : OAI21_X1 port map( B1 => n6076, B2 => n2386, A => n2401, ZN => n3279
                           );
   U2254 : NAND2_X1 port map( A1 => n2386, A2 => n6956, ZN => n2401);
   U2255 : OAI21_X1 port map( B1 => n6075, B2 => n5773, A => n2402, ZN => n3278
                           );
   U2256 : NAND2_X1 port map( A1 => n5773, A2 => n6955, ZN => n2402);
   U2257 : OAI21_X1 port map( B1 => n6074, B2 => n5773, A => n2403, ZN => n3277
                           );
   U2258 : NAND2_X1 port map( A1 => n5773, A2 => n6954, ZN => n2403);
   U2259 : OAI21_X1 port map( B1 => n5499, B2 => n5773, A => n2404, ZN => n3276
                           );
   U2260 : NAND2_X1 port map( A1 => n5774, A2 => n6953, ZN => n2404);
   U2261 : OAI21_X1 port map( B1 => n6072, B2 => n5773, A => n2405, ZN => n3275
                           );
   U2262 : NAND2_X1 port map( A1 => n5774, A2 => n6952, ZN => n2405);
   U2263 : OAI21_X1 port map( B1 => n6071, B2 => n5773, A => n2406, ZN => n3274
                           );
   U2264 : NAND2_X1 port map( A1 => n5774, A2 => n6951, ZN => n2406);
   U2265 : OAI21_X1 port map( B1 => n6070, B2 => n5773, A => n2407, ZN => n3273
                           );
   U2266 : NAND2_X1 port map( A1 => n5774, A2 => n6950, ZN => n2407);
   U2267 : OAI21_X1 port map( B1 => n6069, B2 => n5773, A => n2408, ZN => n3272
                           );
   U2268 : NAND2_X1 port map( A1 => n5774, A2 => n6949, ZN => n2408);
   U2269 : OAI21_X1 port map( B1 => n6068, B2 => n5773, A => n2409, ZN => n3271
                           );
   U2270 : NAND2_X1 port map( A1 => n5774, A2 => n6948, ZN => n2409);
   U2271 : OAI21_X1 port map( B1 => n5481, B2 => n5773, A => n2410, ZN => n3270
                           );
   U2272 : NAND2_X1 port map( A1 => n5774, A2 => n6947, ZN => n2410);
   U2273 : OAI21_X1 port map( B1 => n6066, B2 => n5773, A => n2411, ZN => n3269
                           );
   U2274 : NAND2_X1 port map( A1 => n2386, A2 => n6946, ZN => n2411);
   U2275 : OAI21_X1 port map( B1 => n6065, B2 => n5773, A => n2412, ZN => n3268
                           );
   U2276 : NAND2_X1 port map( A1 => n2386, A2 => n6945, ZN => n2412);
   U2277 : OAI21_X1 port map( B1 => n6064, B2 => n5773, A => n2413, ZN => n3267
                           );
   U2278 : NAND2_X1 port map( A1 => n2386, A2 => n6944, ZN => n2413);
   U2279 : OAI21_X1 port map( B1 => n6063, B2 => n5774, A => n2414, ZN => n3266
                           );
   U2280 : NAND2_X1 port map( A1 => n2386, A2 => n6943, ZN => n2414);
   U2281 : OAI21_X1 port map( B1 => n6062, B2 => n5774, A => n2415, ZN => n3265
                           );
   U2282 : NAND2_X1 port map( A1 => n5774, A2 => n6942, ZN => n2415);
   U2283 : OAI21_X1 port map( B1 => n6061, B2 => n5774, A => n2416, ZN => n3264
                           );
   U2284 : NAND2_X1 port map( A1 => n2386, A2 => n6941, ZN => n2416);
   U2285 : OAI21_X1 port map( B1 => n6060, B2 => n5774, A => n2417, ZN => n3263
                           );
   U2286 : NAND2_X1 port map( A1 => n2386, A2 => n6940, ZN => n2417);
   U2287 : OAI21_X1 port map( B1 => n6059, B2 => n2386, A => n2418, ZN => n3262
                           );
   U2288 : NAND2_X1 port map( A1 => n5773, A2 => n6939, ZN => n2418);
   U2289 : NAND2_X1 port map( A1 => n1555, A2 => n1520, ZN => n2386);
   U2291 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), ZN => n2419);
   U2292 : OAI21_X1 port map( B1 => n6090, B2 => n2420, A => n2421, ZN => n3261
                           );
   U2293 : NAND2_X1 port map( A1 => n609, A2 => n5768, ZN => n2421);
   U2294 : OAI21_X1 port map( B1 => n6089, B2 => n2420, A => n2422, ZN => n3260
                           );
   U2295 : NAND2_X1 port map( A1 => n610, A2 => n5768, ZN => n2422);
   U2296 : OAI21_X1 port map( B1 => n6088, B2 => n2420, A => n2423, ZN => n3259
                           );
   U2297 : NAND2_X1 port map( A1 => n611, A2 => n5768, ZN => n2423);
   U2298 : OAI21_X1 port map( B1 => n6087, B2 => n2420, A => n2424, ZN => n3258
                           );
   U2299 : NAND2_X1 port map( A1 => n612, A2 => n5768, ZN => n2424);
   U2300 : OAI21_X1 port map( B1 => n6086, B2 => n2420, A => n2425, ZN => n3257
                           );
   U2301 : NAND2_X1 port map( A1 => n613, A2 => n5764, ZN => n2425);
   U2302 : OAI21_X1 port map( B1 => n6085, B2 => n2420, A => n2426, ZN => n3256
                           );
   U2303 : NAND2_X1 port map( A1 => n614, A2 => n5764, ZN => n2426);
   U2304 : OAI21_X1 port map( B1 => n6084, B2 => n2420, A => n2427, ZN => n3255
                           );
   U2305 : NAND2_X1 port map( A1 => n615, A2 => n5764, ZN => n2427);
   U2306 : OAI21_X1 port map( B1 => n6083, B2 => n2420, A => n2428, ZN => n3254
                           );
   U2307 : NAND2_X1 port map( A1 => n616, A2 => n2420, ZN => n2428);
   U2308 : OAI21_X1 port map( B1 => n6082, B2 => n2420, A => n2429, ZN => n3253
                           );
   U2309 : NAND2_X1 port map( A1 => n617, A2 => n2420, ZN => n2429);
   U2310 : OAI21_X1 port map( B1 => n5523, B2 => n2420, A => n2430, ZN => n3252
                           );
   U2311 : NAND2_X1 port map( A1 => n618, A2 => n2420, ZN => n2430);
   U2312 : OAI21_X1 port map( B1 => n6080, B2 => n2420, A => n2431, ZN => n3251
                           );
   U2313 : NAND2_X1 port map( A1 => n619, A2 => n2420, ZN => n2431);
   U2314 : OAI21_X1 port map( B1 => n6079, B2 => n2420, A => n2432, ZN => n3250
                           );
   U2315 : NAND2_X1 port map( A1 => n620, A2 => n2420, ZN => n2432);
   U2316 : OAI21_X1 port map( B1 => n6078, B2 => n2420, A => n2433, ZN => n3249
                           );
   U2317 : NAND2_X1 port map( A1 => n621, A2 => n5768, ZN => n2433);
   U2318 : OAI21_X1 port map( B1 => n6077, B2 => n2420, A => n2434, ZN => n3248
                           );
   U2319 : NAND2_X1 port map( A1 => n622, A2 => n5764, ZN => n2434);
   U2320 : OAI21_X1 port map( B1 => n6076, B2 => n2420, A => n2435, ZN => n3247
                           );
   U2321 : NAND2_X1 port map( A1 => n623, A2 => n2420, ZN => n2435);
   U2322 : OAI21_X1 port map( B1 => n6075, B2 => n5768, A => n2436, ZN => n3246
                           );
   U2323 : NAND2_X1 port map( A1 => n624, A2 => n2420, ZN => n2436);
   U2324 : OAI21_X1 port map( B1 => n6074, B2 => n5764, A => n2437, ZN => n3245
                           );
   U2325 : NAND2_X1 port map( A1 => n625, A2 => n5764, ZN => n2437);
   U2326 : OAI21_X1 port map( B1 => n5499, B2 => n5768, A => n2438, ZN => n3244
                           );
   U2327 : NAND2_X1 port map( A1 => n626, A2 => n5764, ZN => n2438);
   U2328 : OAI21_X1 port map( B1 => n6072, B2 => n5764, A => n2439, ZN => n3243
                           );
   U2329 : NAND2_X1 port map( A1 => n627, A2 => n5764, ZN => n2439);
   U2330 : OAI21_X1 port map( B1 => n6071, B2 => n5768, A => n2440, ZN => n3242
                           );
   U2331 : NAND2_X1 port map( A1 => n628, A2 => n5764, ZN => n2440);
   U2332 : OAI21_X1 port map( B1 => n6070, B2 => n5764, A => n2441, ZN => n3241
                           );
   U2333 : NAND2_X1 port map( A1 => n629, A2 => n5764, ZN => n2441);
   U2334 : OAI21_X1 port map( B1 => n6069, B2 => n5768, A => n2442, ZN => n3240
                           );
   U2335 : NAND2_X1 port map( A1 => n630, A2 => n5764, ZN => n2442);
   U2336 : OAI21_X1 port map( B1 => n6068, B2 => n5764, A => n2443, ZN => n3239
                           );
   U2337 : NAND2_X1 port map( A1 => n631, A2 => n5764, ZN => n2443);
   U2338 : OAI21_X1 port map( B1 => n5481, B2 => n5768, A => n2444, ZN => n3238
                           );
   U2339 : NAND2_X1 port map( A1 => n632, A2 => n5764, ZN => n2444);
   U2340 : OAI21_X1 port map( B1 => n6066, B2 => n5764, A => n2445, ZN => n3237
                           );
   U2341 : NAND2_X1 port map( A1 => n633, A2 => n5768, ZN => n2445);
   U2342 : OAI21_X1 port map( B1 => n6065, B2 => n5768, A => n2446, ZN => n3236
                           );
   U2343 : NAND2_X1 port map( A1 => n634, A2 => n5768, ZN => n2446);
   U2344 : OAI21_X1 port map( B1 => n6064, B2 => n5764, A => n2447, ZN => n3235
                           );
   U2345 : NAND2_X1 port map( A1 => n635, A2 => n5768, ZN => n2447);
   U2346 : OAI21_X1 port map( B1 => n6063, B2 => n5768, A => n2448, ZN => n3234
                           );
   U2347 : NAND2_X1 port map( A1 => n636, A2 => n5768, ZN => n2448);
   U2348 : OAI21_X1 port map( B1 => n6062, B2 => n5768, A => n2449, ZN => n3233
                           );
   U2349 : NAND2_X1 port map( A1 => n637, A2 => n5764, ZN => n2449);
   U2350 : OAI21_X1 port map( B1 => n6061, B2 => n5768, A => n2450, ZN => n3232
                           );
   U2351 : NAND2_X1 port map( A1 => n638, A2 => n5764, ZN => n2450);
   U2352 : OAI21_X1 port map( B1 => n6060, B2 => n5768, A => n2451, ZN => n3231
                           );
   U2353 : NAND2_X1 port map( A1 => n639, A2 => n2420, ZN => n2451);
   U2354 : OAI21_X1 port map( B1 => n6059, B2 => n2420, A => n2452, ZN => n3230
                           );
   U2355 : NAND2_X1 port map( A1 => n640, A2 => n5768, ZN => n2452);
   U2356 : NAND2_X1 port map( A1 => n1778, A2 => n1520, ZN => n2420);
   U2357 : NOR2_X1 port map( A1 => n2453, A2 => n6050, ZN => n1778);
   U2358 : NAND2_X1 port map( A1 => n2454, A2 => n2455, ZN => n3229);
   U2359 : NOR4_X1 port map( A1 => n2456, A2 => n2457, A3 => n2458, A4 => n2459
                           , ZN => n2455);
   U2360 : OAI21_X1 port map( B1 => n1423, B2 => n5762, A => n2461, ZN => n2459
                           );
   U2361 : NAND2_X1 port map( A1 => n5759, A2 => n6859, ZN => n2461);
   U2362 : OAI21_X1 port map( B1 => n6059, B2 => n5756, A => n2464, ZN => n2458
                           );
   U2363 : AOI22_X1 port map( A1 => n5753, A2 => n6707, B1 => n5750, B2 => 
                           n6987, ZN => n2464);
   U2364 : NAND2_X1 port map( A1 => n2467, A2 => n2468, ZN => n2457);
   U2365 : AOI22_X1 port map( A1 => n5745, A2 => n2830, B1 => n5744, B2 => 
                           n6938, ZN => n2468);
   U2366 : AOI22_X1 port map( A1 => n5741, A2 => n6604, B1 => n5738, B2 => 
                           n7051, ZN => n2467);
   U2368 : AOI22_X1 port map( A1 => n5735, A2 => n6742, B1 => n5732, B2 => 
                           n7019, ZN => n2476);
   U2369 : AOI22_X1 port map( A1 => n5729, A2 => n6667, B1 => n2480, B2 => 
                           n6937, ZN => n2475);
   U2370 : AOI22_X1 port map( A1 => n5723, A2 => n6710, B1 => n5720, B2 => 
                           n2382, ZN => n2474);
   U2371 : AOI22_X1 port map( A1 => n5717, A2 => n640, B1 => n5714, B2 => n480,
                           ZN => n2473);
   U2372 : NOR4_X1 port map( A1 => n2485, A2 => n2486, A3 => n2487, A4 => n2488
                           , ZN => n2454);
   U2373 : NAND2_X1 port map( A1 => n2489, A2 => n2490, ZN => n2488);
   U2374 : AOI22_X1 port map( A1 => n5711, A2 => n416, B1 => n5708, B2 => n7083
                           , ZN => n2490);
   U2375 : AOI22_X1 port map( A1 => n5705, A2 => n6796, B1 => n5934, B2 => 
                           OUT1_31_port, ZN => n2489);
   U2376 : NAND2_X1 port map( A1 => n2494, A2 => n2495, ZN => n2487);
   U2377 : AOI22_X1 port map( A1 => n2496, A2 => n448, B1 => n5697, B2 => n6939
                           , ZN => n2495);
   U2378 : AOI22_X1 port map( A1 => n5696, A2 => n6764, B1 => n5693, B2 => n576
                           , ZN => n2494);
   U2379 : NAND2_X1 port map( A1 => n2500, A2 => n2501, ZN => n2486);
   U2380 : AOI22_X1 port map( A1 => n5690, A2 => n704, B1 => n5687, B2 => n672,
                           ZN => n2501);
   U2381 : AOI22_X1 port map( A1 => n5684, A2 => n736, B1 => n5681, B2 => n608,
                           ZN => n2500);
   U2382 : NAND2_X1 port map( A1 => n2506, A2 => n2507, ZN => n2485);
   U2383 : AOI22_X1 port map( A1 => n2508, A2 => n512, B1 => n5673, B2 => n384,
                           ZN => n2507);
   U2384 : AOI22_X1 port map( A1 => n5672, A2 => n544, B1 => n5669, B2 => n352,
                           ZN => n2506);
   U2385 : NAND2_X1 port map( A1 => n2512, A2 => n2513, ZN => n3228);
   U2386 : NOR4_X1 port map( A1 => n2514, A2 => n2515, A3 => n2516, A4 => n2517
                           , ZN => n2513);
   U2387 : OAI21_X1 port map( B1 => n1424, B2 => n5762, A => n2518, ZN => n2517
                           );
   U2388 : NAND2_X1 port map( A1 => n5759, A2 => n6858, ZN => n2518);
   U2389 : OAI21_X1 port map( B1 => n6060, B2 => n5756, A => n2519, ZN => n2516
                           );
   U2390 : AOI22_X1 port map( A1 => n5753, A2 => n6706, B1 => n5750, B2 => 
                           n6986, ZN => n2519);
   U2391 : NAND2_X1 port map( A1 => n2520, A2 => n2521, ZN => n2515);
   U2392 : AOI22_X1 port map( A1 => n5745, A2 => n2829, B1 => n5744, B2 => 
                           n6936, ZN => n2521);
   U2393 : AOI22_X1 port map( A1 => n5741, A2 => n6605, B1 => n5738, B2 => 
                           n7050, ZN => n2520);
   U2395 : AOI22_X1 port map( A1 => n5735, A2 => n6741, B1 => n5732, B2 => 
                           n7018, ZN => n2525);
   U2396 : AOI22_X1 port map( A1 => n5729, A2 => n6666, B1 => n2480, B2 => 
                           n6935, ZN => n2524);
   U2397 : AOI22_X1 port map( A1 => n5723, A2 => n6709, B1 => n5720, B2 => 
                           n2379, ZN => n2523);
   U2398 : AOI22_X1 port map( A1 => n5717, A2 => n639, B1 => n5714, B2 => n479,
                           ZN => n2522);
   U2399 : NOR4_X1 port map( A1 => n2526, A2 => n2527, A3 => n2528, A4 => n2529
                           , ZN => n2512);
   U2400 : NAND2_X1 port map( A1 => n2530, A2 => n2531, ZN => n2529);
   U2401 : AOI22_X1 port map( A1 => n5711, A2 => n415, B1 => n5708, B2 => n7082
                           , ZN => n2531);
   U2402 : AOI22_X1 port map( A1 => n5705, A2 => n6797, B1 => n5934, B2 => 
                           OUT1_30_port, ZN => n2530);
   U2403 : NAND2_X1 port map( A1 => n2532, A2 => n2533, ZN => n2528);
   U2404 : AOI22_X1 port map( A1 => n2496, A2 => n447, B1 => n5697, B2 => n6940
                           , ZN => n2533);
   U2405 : AOI22_X1 port map( A1 => n5696, A2 => n6765, B1 => n5693, B2 => n575
                           , ZN => n2532);
   U2406 : NAND2_X1 port map( A1 => n2534, A2 => n2535, ZN => n2527);
   U2407 : AOI22_X1 port map( A1 => n5690, A2 => n703, B1 => n5687, B2 => n671,
                           ZN => n2535);
   U2408 : AOI22_X1 port map( A1 => n5684, A2 => n735, B1 => n5681, B2 => n607,
                           ZN => n2534);
   U2409 : NAND2_X1 port map( A1 => n2536, A2 => n2537, ZN => n2526);
   U2410 : AOI22_X1 port map( A1 => n2508, A2 => n511, B1 => n5673, B2 => n383,
                           ZN => n2537);
   U2411 : AOI22_X1 port map( A1 => n5672, A2 => n543, B1 => n5669, B2 => n351,
                           ZN => n2536);
   U2412 : NAND2_X1 port map( A1 => n2538, A2 => n2539, ZN => n3227);
   U2413 : NOR4_X1 port map( A1 => n2540, A2 => n2541, A3 => n2542, A4 => n2543
                           , ZN => n2539);
   U2414 : OAI21_X1 port map( B1 => n1425, B2 => n5762, A => n2544, ZN => n2543
                           );
   U2415 : NAND2_X1 port map( A1 => n5759, A2 => n6857, ZN => n2544);
   U2416 : OAI21_X1 port map( B1 => n6061, B2 => n5756, A => n2545, ZN => n2542
                           );
   U2417 : AOI22_X1 port map( A1 => n5753, A2 => n6705, B1 => n5750, B2 => 
                           n6985, ZN => n2545);
   U2418 : NAND2_X1 port map( A1 => n2546, A2 => n2547, ZN => n2541);
   U2419 : AOI22_X1 port map( A1 => n5745, A2 => n2828, B1 => n5744, B2 => 
                           n6934, ZN => n2547);
   U2420 : AOI22_X1 port map( A1 => n5741, A2 => n6606, B1 => n5738, B2 => 
                           n7049, ZN => n2546);
   U2422 : AOI22_X1 port map( A1 => n5735, A2 => n6740, B1 => n5732, B2 => 
                           n7017, ZN => n2551);
   U2423 : AOI22_X1 port map( A1 => n5729, A2 => n6665, B1 => n2480, B2 => 
                           n6933, ZN => n2550);
   U2424 : AOI22_X1 port map( A1 => n5723, A2 => n6708, B1 => n5720, B2 => 
                           n2376, ZN => n2549);
   U2425 : AOI22_X1 port map( A1 => n5717, A2 => n638, B1 => n5714, B2 => n478,
                           ZN => n2548);
   U2426 : NOR4_X1 port map( A1 => n2552, A2 => n2553, A3 => n2554, A4 => n2555
                           , ZN => n2538);
   U2427 : NAND2_X1 port map( A1 => n2556, A2 => n2557, ZN => n2555);
   U2428 : AOI22_X1 port map( A1 => n5711, A2 => n414, B1 => n5708, B2 => n7081
                           , ZN => n2557);
   U2429 : AOI22_X1 port map( A1 => n5705, A2 => n6798, B1 => n5935, B2 => 
                           OUT1_29_port, ZN => n2556);
   U2430 : NAND2_X1 port map( A1 => n2558, A2 => n2559, ZN => n2554);
   U2431 : AOI22_X1 port map( A1 => n2496, A2 => n446, B1 => n5697, B2 => n6941
                           , ZN => n2559);
   U2432 : AOI22_X1 port map( A1 => n5696, A2 => n6766, B1 => n5693, B2 => n574
                           , ZN => n2558);
   U2433 : NAND2_X1 port map( A1 => n2560, A2 => n2561, ZN => n2553);
   U2434 : AOI22_X1 port map( A1 => n5690, A2 => n702, B1 => n5687, B2 => n670,
                           ZN => n2561);
   U2435 : AOI22_X1 port map( A1 => n5684, A2 => n734, B1 => n5681, B2 => n606,
                           ZN => n2560);
   U2436 : NAND2_X1 port map( A1 => n2562, A2 => n2563, ZN => n2552);
   U2437 : AOI22_X1 port map( A1 => n2508, A2 => n510, B1 => n5673, B2 => n382,
                           ZN => n2563);
   U2438 : AOI22_X1 port map( A1 => n5672, A2 => n542, B1 => n5669, B2 => n350,
                           ZN => n2562);
   U2439 : NAND2_X1 port map( A1 => n2564, A2 => n2565, ZN => n3226);
   U2440 : NOR4_X1 port map( A1 => n2566, A2 => n2567, A3 => n2568, A4 => n2569
                           , ZN => n2565);
   U2441 : OAI21_X1 port map( B1 => n1426, B2 => n5762, A => n2570, ZN => n2569
                           );
   U2442 : NAND2_X1 port map( A1 => n5759, A2 => n6856, ZN => n2570);
   U2443 : OAI21_X1 port map( B1 => n6062, B2 => n5756, A => n2571, ZN => n2568
                           );
   U2444 : AOI22_X1 port map( A1 => n5753, A2 => n6704, B1 => n5750, B2 => 
                           n6984, ZN => n2571);
   U2445 : NAND2_X1 port map( A1 => n2572, A2 => n2573, ZN => n2567);
   U2446 : AOI22_X1 port map( A1 => n5745, A2 => n2827, B1 => n5744, B2 => 
                           n6932, ZN => n2573);
   U2447 : AOI22_X1 port map( A1 => n5741, A2 => n6607, B1 => n5738, B2 => 
                           n7048, ZN => n2572);
   U2449 : AOI22_X1 port map( A1 => n5735, A2 => n6739, B1 => n5732, B2 => 
                           n7016, ZN => n2577);
   U2450 : AOI22_X1 port map( A1 => n5729, A2 => n6664, B1 => n2480, B2 => 
                           n6931, ZN => n2576);
   U2451 : AOI22_X1 port map( A1 => n5723, A2 => n2270, B1 => n5720, B2 => 
                           n2373, ZN => n2575);
   U2452 : AOI22_X1 port map( A1 => n5717, A2 => n637, B1 => n5714, B2 => n477,
                           ZN => n2574);
   U2453 : NOR4_X1 port map( A1 => n2578, A2 => n2579, A3 => n2580, A4 => n2581
                           , ZN => n2564);
   U2454 : NAND2_X1 port map( A1 => n2582, A2 => n2583, ZN => n2581);
   U2455 : AOI22_X1 port map( A1 => n5711, A2 => n413, B1 => n5708, B2 => n7080
                           , ZN => n2583);
   U2456 : AOI22_X1 port map( A1 => n5705, A2 => n6799, B1 => n5932, B2 => 
                           OUT1_28_port, ZN => n2582);
   U2457 : NAND2_X1 port map( A1 => n2584, A2 => n2585, ZN => n2580);
   U2458 : AOI22_X1 port map( A1 => n2496, A2 => n445, B1 => n5697, B2 => n6942
                           , ZN => n2585);
   U2459 : AOI22_X1 port map( A1 => n5696, A2 => n6767, B1 => n5693, B2 => n573
                           , ZN => n2584);
   U2460 : NAND2_X1 port map( A1 => n2586, A2 => n2587, ZN => n2579);
   U2461 : AOI22_X1 port map( A1 => n5690, A2 => n701, B1 => n5687, B2 => n669,
                           ZN => n2587);
   U2462 : AOI22_X1 port map( A1 => n5684, A2 => n733, B1 => n5681, B2 => n605,
                           ZN => n2586);
   U2463 : NAND2_X1 port map( A1 => n2588, A2 => n2589, ZN => n2578);
   U2464 : AOI22_X1 port map( A1 => n2508, A2 => n509, B1 => n5673, B2 => n381,
                           ZN => n2589);
   U2465 : AOI22_X1 port map( A1 => n5672, A2 => n541, B1 => n5669, B2 => n349,
                           ZN => n2588);
   U2466 : NAND2_X1 port map( A1 => n2590, A2 => n2591, ZN => n3225);
   U2467 : NOR4_X1 port map( A1 => n2592, A2 => n2593, A3 => n2594, A4 => n2595
                           , ZN => n2591);
   U2468 : OAI21_X1 port map( B1 => n1427, B2 => n5762, A => n2596, ZN => n2595
                           );
   U2469 : NAND2_X1 port map( A1 => n5759, A2 => n6855, ZN => n2596);
   U2470 : OAI21_X1 port map( B1 => n6063, B2 => n5756, A => n2597, ZN => n2594
                           );
   U2471 : AOI22_X1 port map( A1 => n5753, A2 => n6703, B1 => n5750, B2 => 
                           n6983, ZN => n2597);
   U2472 : NAND2_X1 port map( A1 => n2598, A2 => n2599, ZN => n2593);
   U2473 : AOI22_X1 port map( A1 => n5745, A2 => n2826, B1 => n5744, B2 => 
                           n6930, ZN => n2599);
   U2474 : AOI22_X1 port map( A1 => n5741, A2 => n6608, B1 => n5738, B2 => 
                           n7047, ZN => n2598);
   U2476 : AOI22_X1 port map( A1 => n5735, A2 => n6738, B1 => n5732, B2 => 
                           n7015, ZN => n2603);
   U2477 : AOI22_X1 port map( A1 => n5729, A2 => n6663, B1 => n2480, B2 => 
                           n6929, ZN => n2602);
   U2478 : AOI22_X1 port map( A1 => n5723, A2 => n2265, B1 => n5720, B2 => 
                           n2370, ZN => n2601);
   U2479 : AOI22_X1 port map( A1 => n5717, A2 => n636, B1 => n5714, B2 => n476,
                           ZN => n2600);
   U2480 : NOR4_X1 port map( A1 => n2604, A2 => n2605, A3 => n2606, A4 => n2607
                           , ZN => n2590);
   U2481 : NAND2_X1 port map( A1 => n2608, A2 => n2609, ZN => n2607);
   U2482 : AOI22_X1 port map( A1 => n5711, A2 => n412, B1 => n5708, B2 => n7079
                           , ZN => n2609);
   U2483 : AOI22_X1 port map( A1 => n5705, A2 => n6800, B1 => n5935, B2 => 
                           OUT1_27_port, ZN => n2608);
   U2484 : NAND2_X1 port map( A1 => n2610, A2 => n2611, ZN => n2606);
   U2485 : AOI22_X1 port map( A1 => n5701, A2 => n444, B1 => n5697, B2 => n6943
                           , ZN => n2611);
   U2486 : AOI22_X1 port map( A1 => n5696, A2 => n6768, B1 => n5693, B2 => n572
                           , ZN => n2610);
   U2487 : NAND2_X1 port map( A1 => n2612, A2 => n2613, ZN => n2605);
   U2488 : AOI22_X1 port map( A1 => n5690, A2 => n700, B1 => n5687, B2 => n668,
                           ZN => n2613);
   U2489 : AOI22_X1 port map( A1 => n5684, A2 => n732, B1 => n5681, B2 => n604,
                           ZN => n2612);
   U2490 : NAND2_X1 port map( A1 => n2614, A2 => n2615, ZN => n2604);
   U2491 : AOI22_X1 port map( A1 => n5677, A2 => n508, B1 => n5673, B2 => n380,
                           ZN => n2615);
   U2492 : AOI22_X1 port map( A1 => n5672, A2 => n540, B1 => n5669, B2 => n348,
                           ZN => n2614);
   U2493 : NAND2_X1 port map( A1 => n2616, A2 => n2617, ZN => n3224);
   U2494 : NOR4_X1 port map( A1 => n2618, A2 => n2619, A3 => n2620, A4 => n2621
                           , ZN => n2617);
   U2495 : OAI21_X1 port map( B1 => n1428, B2 => n5762, A => n2622, ZN => n2621
                           );
   U2496 : NAND2_X1 port map( A1 => n5759, A2 => n6854, ZN => n2622);
   U2497 : OAI21_X1 port map( B1 => n6064, B2 => n5756, A => n2623, ZN => n2620
                           );
   U2498 : AOI22_X1 port map( A1 => n5753, A2 => n6702, B1 => n5750, B2 => 
                           n6982, ZN => n2623);
   U2499 : NAND2_X1 port map( A1 => n2624, A2 => n2625, ZN => n2619);
   U2500 : AOI22_X1 port map( A1 => n5745, A2 => n2825, B1 => n5744, B2 => 
                           n6928, ZN => n2625);
   U2501 : AOI22_X1 port map( A1 => n5741, A2 => n6609, B1 => n5738, B2 => 
                           n7046, ZN => n2624);
   U2503 : AOI22_X1 port map( A1 => n5735, A2 => n6737, B1 => n5732, B2 => 
                           n7014, ZN => n2629);
   U2504 : AOI22_X1 port map( A1 => n5729, A2 => n6662, B1 => n2480, B2 => 
                           n6927, ZN => n2628);
   U2505 : AOI22_X1 port map( A1 => n5723, A2 => n2260, B1 => n5720, B2 => 
                           n2367, ZN => n2627);
   U2506 : AOI22_X1 port map( A1 => n5717, A2 => n635, B1 => n5714, B2 => n475,
                           ZN => n2626);
   U2507 : NOR4_X1 port map( A1 => n2630, A2 => n2631, A3 => n2632, A4 => n2633
                           , ZN => n2616);
   U2508 : NAND2_X1 port map( A1 => n2634, A2 => n2635, ZN => n2633);
   U2509 : AOI22_X1 port map( A1 => n5711, A2 => n411, B1 => n5708, B2 => n7078
                           , ZN => n2635);
   U2510 : AOI22_X1 port map( A1 => n5705, A2 => n6801, B1 => n5934, B2 => 
                           OUT1_26_port, ZN => n2634);
   U2511 : NAND2_X1 port map( A1 => n2636, A2 => n2637, ZN => n2632);
   U2512 : AOI22_X1 port map( A1 => n5701, A2 => n443, B1 => n5697, B2 => n6944
                           , ZN => n2637);
   U2513 : AOI22_X1 port map( A1 => n5696, A2 => n6769, B1 => n5693, B2 => n571
                           , ZN => n2636);
   U2514 : NAND2_X1 port map( A1 => n2638, A2 => n2639, ZN => n2631);
   U2515 : AOI22_X1 port map( A1 => n5690, A2 => n699, B1 => n5687, B2 => n667,
                           ZN => n2639);
   U2516 : AOI22_X1 port map( A1 => n5684, A2 => n731, B1 => n5681, B2 => n603,
                           ZN => n2638);
   U2517 : NAND2_X1 port map( A1 => n2640, A2 => n2641, ZN => n2630);
   U2518 : AOI22_X1 port map( A1 => n5677, A2 => n507, B1 => n5673, B2 => n379,
                           ZN => n2641);
   U2519 : AOI22_X1 port map( A1 => n5672, A2 => n539, B1 => n5669, B2 => n347,
                           ZN => n2640);
   U2520 : NAND2_X1 port map( A1 => n2642, A2 => n2643, ZN => n3223);
   U2521 : NOR4_X1 port map( A1 => n2644, A2 => n2645, A3 => n2646, A4 => n2647
                           , ZN => n2643);
   U2522 : OAI21_X1 port map( B1 => n1429, B2 => n5762, A => n2648, ZN => n2647
                           );
   U2523 : NAND2_X1 port map( A1 => n5759, A2 => n6853, ZN => n2648);
   U2524 : OAI21_X1 port map( B1 => n6065, B2 => n5756, A => n2649, ZN => n2646
                           );
   U2525 : AOI22_X1 port map( A1 => n5753, A2 => n6701, B1 => n5750, B2 => 
                           n6981, ZN => n2649);
   U2526 : NAND2_X1 port map( A1 => n2650, A2 => n2651, ZN => n2645);
   U2527 : AOI22_X1 port map( A1 => n5745, A2 => n2824, B1 => n5744, B2 => 
                           n6926, ZN => n2651);
   U2528 : AOI22_X1 port map( A1 => n5741, A2 => n6610, B1 => n5738, B2 => 
                           n7045, ZN => n2650);
   U2530 : AOI22_X1 port map( A1 => n5735, A2 => n6736, B1 => n5732, B2 => 
                           n7013, ZN => n2655);
   U2531 : AOI22_X1 port map( A1 => n5729, A2 => n6661, B1 => n2480, B2 => 
                           n6925, ZN => n2654);
   U2532 : AOI22_X1 port map( A1 => n5723, A2 => n2255, B1 => n5720, B2 => 
                           n2364, ZN => n2653);
   U2533 : AOI22_X1 port map( A1 => n5717, A2 => n634, B1 => n5714, B2 => n474,
                           ZN => n2652);
   U2534 : NOR4_X1 port map( A1 => n2656, A2 => n2657, A3 => n2658, A4 => n2659
                           , ZN => n2642);
   U2535 : NAND2_X1 port map( A1 => n2660, A2 => n2661, ZN => n2659);
   U2536 : AOI22_X1 port map( A1 => n5711, A2 => n410, B1 => n5708, B2 => n7077
                           , ZN => n2661);
   U2537 : AOI22_X1 port map( A1 => n5705, A2 => n6802, B1 => n5935, B2 => 
                           OUT1_25_port, ZN => n2660);
   U2538 : NAND2_X1 port map( A1 => n2662, A2 => n2663, ZN => n2658);
   U2539 : AOI22_X1 port map( A1 => n2496, A2 => n442, B1 => n2497, B2 => n6945
                           , ZN => n2663);
   U2540 : AOI22_X1 port map( A1 => n5696, A2 => n6770, B1 => n5693, B2 => n570
                           , ZN => n2662);
   U2541 : NAND2_X1 port map( A1 => n2664, A2 => n2665, ZN => n2657);
   U2542 : AOI22_X1 port map( A1 => n5690, A2 => n698, B1 => n5687, B2 => n666,
                           ZN => n2665);
   U2543 : AOI22_X1 port map( A1 => n5684, A2 => n730, B1 => n5681, B2 => n602,
                           ZN => n2664);
   U2544 : NAND2_X1 port map( A1 => n2666, A2 => n2667, ZN => n2656);
   U2545 : AOI22_X1 port map( A1 => n2508, A2 => n506, B1 => n2509, B2 => n378,
                           ZN => n2667);
   U2546 : AOI22_X1 port map( A1 => n5672, A2 => n538, B1 => n5669, B2 => n346,
                           ZN => n2666);
   U2547 : NAND2_X1 port map( A1 => n2668, A2 => n2669, ZN => n3222);
   U2548 : NOR4_X1 port map( A1 => n2670, A2 => n2671, A3 => n2672, A4 => n2673
                           , ZN => n2669);
   U2549 : OAI21_X1 port map( B1 => n1430, B2 => n5762, A => n2674, ZN => n2673
                           );
   U2550 : NAND2_X1 port map( A1 => n5759, A2 => n6852, ZN => n2674);
   U2551 : OAI21_X1 port map( B1 => n6066, B2 => n5756, A => n2675, ZN => n2672
                           );
   U2552 : AOI22_X1 port map( A1 => n5753, A2 => n6700, B1 => n5750, B2 => 
                           n6980, ZN => n2675);
   U2553 : NAND2_X1 port map( A1 => n2676, A2 => n2677, ZN => n2671);
   U2554 : AOI22_X1 port map( A1 => n2469, A2 => n2823, B1 => n5744, B2 => 
                           n6924, ZN => n2677);
   U2555 : AOI22_X1 port map( A1 => n5741, A2 => n6611, B1 => n5738, B2 => 
                           n7044, ZN => n2676);
   U2557 : AOI22_X1 port map( A1 => n5735, A2 => n6735, B1 => n5732, B2 => 
                           n7012, ZN => n2681);
   U2558 : AOI22_X1 port map( A1 => n5729, A2 => n6660, B1 => n5725, B2 => 
                           n6923, ZN => n2680);
   U2559 : AOI22_X1 port map( A1 => n5723, A2 => n2250, B1 => n5720, B2 => 
                           n2361, ZN => n2679);
   U2560 : AOI22_X1 port map( A1 => n5717, A2 => n633, B1 => n5714, B2 => n473,
                           ZN => n2678);
   U2561 : NOR4_X1 port map( A1 => n2682, A2 => n2683, A3 => n2684, A4 => n2685
                           , ZN => n2668);
   U2562 : NAND2_X1 port map( A1 => n2686, A2 => n2687, ZN => n2685);
   U2563 : AOI22_X1 port map( A1 => n5711, A2 => n409, B1 => n5708, B2 => n7076
                           , ZN => n2687);
   U2564 : AOI22_X1 port map( A1 => n5705, A2 => n6803, B1 => n5935, B2 => 
                           OUT1_24_port, ZN => n2686);
   U2565 : NAND2_X1 port map( A1 => n2688, A2 => n2689, ZN => n2684);
   U2566 : AOI22_X1 port map( A1 => n2496, A2 => n441, B1 => n2497, B2 => n6946
                           , ZN => n2689);
   U2567 : AOI22_X1 port map( A1 => n5696, A2 => n6771, B1 => n5693, B2 => n569
                           , ZN => n2688);
   U2568 : NAND2_X1 port map( A1 => n2690, A2 => n2691, ZN => n2683);
   U2569 : AOI22_X1 port map( A1 => n5690, A2 => n697, B1 => n5687, B2 => n665,
                           ZN => n2691);
   U2570 : AOI22_X1 port map( A1 => n5684, A2 => n729, B1 => n5681, B2 => n601,
                           ZN => n2690);
   U2571 : NAND2_X1 port map( A1 => n2692, A2 => n2693, ZN => n2682);
   U2572 : AOI22_X1 port map( A1 => n2508, A2 => n505, B1 => n2509, B2 => n377,
                           ZN => n2693);
   U2573 : AOI22_X1 port map( A1 => n5672, A2 => n537, B1 => n5669, B2 => n345,
                           ZN => n2692);
   U2574 : NAND2_X1 port map( A1 => n2694, A2 => n2695, ZN => n3221);
   U2575 : NOR4_X1 port map( A1 => n2696, A2 => n2697, A3 => n2698, A4 => n2699
                           , ZN => n2695);
   U2576 : OAI21_X1 port map( B1 => n1431, B2 => n2460, A => n2700, ZN => n2699
                           );
   U2577 : NAND2_X1 port map( A1 => n5759, A2 => n6851, ZN => n2700);
   U2578 : OAI21_X1 port map( B1 => n5481, B2 => n2463, A => n2701, ZN => n2698
                           );
   U2579 : AOI22_X1 port map( A1 => n5753, A2 => n6699, B1 => n2466, B2 => 
                           n6979, ZN => n2701);
   U2580 : NAND2_X1 port map( A1 => n2702, A2 => n2703, ZN => n2697);
   U2581 : AOI22_X1 port map( A1 => n5745, A2 => n2822, B1 => n2470, B2 => 
                           n6922, ZN => n2703);
   U2582 : AOI22_X1 port map( A1 => n2471, A2 => n6612, B1 => n5738, B2 => 
                           n7043, ZN => n2702);
   U2584 : AOI22_X1 port map( A1 => n5735, A2 => n6734, B1 => n2478, B2 => 
                           n7011, ZN => n2707);
   U2585 : AOI22_X1 port map( A1 => n5729, A2 => n6659, B1 => n5725, B2 => 
                           n6921, ZN => n2706);
   U2586 : AOI22_X1 port map( A1 => n2481, A2 => n2245, B1 => n5720, B2 => 
                           n2358, ZN => n2705);
   U2587 : AOI22_X1 port map( A1 => n2483, A2 => n632, B1 => n5714, B2 => n472,
                           ZN => n2704);
   U2588 : NOR4_X1 port map( A1 => n2708, A2 => n2709, A3 => n2710, A4 => n2711
                           , ZN => n2694);
   U2589 : NAND2_X1 port map( A1 => n2712, A2 => n2713, ZN => n2711);
   U2590 : AOI22_X1 port map( A1 => n2491, A2 => n408, B1 => n5708, B2 => n7075
                           , ZN => n2713);
   U2591 : AOI22_X1 port map( A1 => n5705, A2 => n6804, B1 => n5935, B2 => 
                           OUT1_23_port, ZN => n2712);
   U2592 : NAND2_X1 port map( A1 => n2714, A2 => n2715, ZN => n2710);
   U2593 : AOI22_X1 port map( A1 => n5701, A2 => n440, B1 => n2497, B2 => n6947
                           , ZN => n2715);
   U2594 : AOI22_X1 port map( A1 => n5696, A2 => n6772, B1 => n2499, B2 => n568
                           , ZN => n2714);
   U2595 : NAND2_X1 port map( A1 => n2716, A2 => n2717, ZN => n2709);
   U2596 : AOI22_X1 port map( A1 => n5690, A2 => n696, B1 => n2503, B2 => n664,
                           ZN => n2717);
   U2597 : AOI22_X1 port map( A1 => n5684, A2 => n728, B1 => n2505, B2 => n600,
                           ZN => n2716);
   U2598 : NAND2_X1 port map( A1 => n2718, A2 => n2719, ZN => n2708);
   U2599 : AOI22_X1 port map( A1 => n5677, A2 => n504, B1 => n2509, B2 => n376,
                           ZN => n2719);
   U2600 : AOI22_X1 port map( A1 => n5672, A2 => n536, B1 => n2511, B2 => n344,
                           ZN => n2718);
   U2601 : NAND2_X1 port map( A1 => n2720, A2 => n2721, ZN => n3220);
   U2602 : NOR4_X1 port map( A1 => n2722, A2 => n2723, A3 => n2724, A4 => n2725
                           , ZN => n2721);
   U2603 : OAI21_X1 port map( B1 => n1432, B2 => n2460, A => n2726, ZN => n2725
                           );
   U2604 : NAND2_X1 port map( A1 => n5759, A2 => n6850, ZN => n2726);
   U2605 : OAI21_X1 port map( B1 => n6068, B2 => n2463, A => n2727, ZN => n2724
                           );
   U2606 : AOI22_X1 port map( A1 => n2465, A2 => n6698, B1 => n5750, B2 => 
                           n6978, ZN => n2727);
   U2607 : NAND2_X1 port map( A1 => n2728, A2 => n2729, ZN => n2723);
   U2608 : AOI22_X1 port map( A1 => n2469, A2 => n2821, B1 => n5744, B2 => 
                           n6920, ZN => n2729);
   U2609 : AOI22_X1 port map( A1 => n5741, A2 => n6613, B1 => n2472, B2 => 
                           n7042, ZN => n2728);
   U2611 : AOI22_X1 port map( A1 => n5735, A2 => n6733, B1 => n2478, B2 => 
                           n7010, ZN => n2733);
   U2612 : AOI22_X1 port map( A1 => n5729, A2 => n6658, B1 => n5725, B2 => 
                           n6919, ZN => n2732);
   U2613 : AOI22_X1 port map( A1 => n2481, A2 => n2240, B1 => n5720, B2 => 
                           n2355, ZN => n2731);
   U2614 : AOI22_X1 port map( A1 => n2483, A2 => n631, B1 => n5714, B2 => n471,
                           ZN => n2730);
   U2615 : NOR4_X1 port map( A1 => n2734, A2 => n2735, A3 => n2736, A4 => n2737
                           , ZN => n2720);
   U2616 : NAND2_X1 port map( A1 => n2738, A2 => n2739, ZN => n2737);
   U2617 : AOI22_X1 port map( A1 => n5711, A2 => n407, B1 => n2492, B2 => n7074
                           , ZN => n2739);
   U2618 : AOI22_X1 port map( A1 => n5705, A2 => n6805, B1 => n5935, B2 => 
                           OUT1_22_port, ZN => n2738);
   U2619 : NAND2_X1 port map( A1 => n2740, A2 => n2741, ZN => n2736);
   U2620 : AOI22_X1 port map( A1 => n5701, A2 => n439, B1 => n5697, B2 => n6948
                           , ZN => n2741);
   U2621 : AOI22_X1 port map( A1 => n5696, A2 => n6773, B1 => n2499, B2 => n567
                           , ZN => n2740);
   U2622 : NAND2_X1 port map( A1 => n2742, A2 => n2743, ZN => n2735);
   U2623 : AOI22_X1 port map( A1 => n5690, A2 => n695, B1 => n2503, B2 => n663,
                           ZN => n2743);
   U2624 : AOI22_X1 port map( A1 => n5684, A2 => n727, B1 => n2505, B2 => n599,
                           ZN => n2742);
   U2625 : NAND2_X1 port map( A1 => n2744, A2 => n2745, ZN => n2734);
   U2626 : AOI22_X1 port map( A1 => n5677, A2 => n503, B1 => n5673, B2 => n375,
                           ZN => n2745);
   U2627 : AOI22_X1 port map( A1 => n5672, A2 => n535, B1 => n2511, B2 => n343,
                           ZN => n2744);
   U2628 : NAND2_X1 port map( A1 => n2746, A2 => n2747, ZN => n3219);
   U2629 : NOR4_X1 port map( A1 => n2748, A2 => n2749, A3 => n2750, A4 => n2751
                           , ZN => n2747);
   U2630 : OAI21_X1 port map( B1 => n1433, B2 => n2460, A => n2752, ZN => n2751
                           );
   U2631 : NAND2_X1 port map( A1 => n5759, A2 => n6849, ZN => n2752);
   U2632 : OAI21_X1 port map( B1 => n6069, B2 => n2463, A => n2753, ZN => n2750
                           );
   U2633 : AOI22_X1 port map( A1 => n2465, A2 => n6697, B1 => n5750, B2 => 
                           n6977, ZN => n2753);
   U2634 : NAND2_X1 port map( A1 => n2754, A2 => n2755, ZN => n2749);
   U2635 : AOI22_X1 port map( A1 => n2469, A2 => n2820, B1 => n2470, B2 => 
                           n6918, ZN => n2755);
   U2636 : AOI22_X1 port map( A1 => n5741, A2 => n6614, B1 => n2472, B2 => 
                           n7041, ZN => n2754);
   U2638 : AOI22_X1 port map( A1 => n5735, A2 => n6732, B1 => n2478, B2 => 
                           n7009, ZN => n2759);
   U2639 : AOI22_X1 port map( A1 => n5729, A2 => n6657, B1 => n5725, B2 => 
                           n6917, ZN => n2758);
   U2640 : AOI22_X1 port map( A1 => n2481, A2 => n2235, B1 => n5720, B2 => 
                           n2352, ZN => n2757);
   U2641 : AOI22_X1 port map( A1 => n2483, A2 => n630, B1 => n5714, B2 => n470,
                           ZN => n2756);
   U2642 : NOR4_X1 port map( A1 => n2760, A2 => n2761, A3 => n2762, A4 => n2763
                           , ZN => n2746);
   U2643 : NAND2_X1 port map( A1 => n2764, A2 => n2765, ZN => n2763);
   U2644 : AOI22_X1 port map( A1 => n5711, A2 => n406, B1 => n2492, B2 => n7073
                           , ZN => n2765);
   U2645 : AOI22_X1 port map( A1 => n5705, A2 => n6806, B1 => n5935, B2 => 
                           OUT1_21_port, ZN => n2764);
   U2646 : NAND2_X1 port map( A1 => n2766, A2 => n2767, ZN => n2762);
   U2647 : AOI22_X1 port map( A1 => n5701, A2 => n438, B1 => n2497, B2 => n6949
                           , ZN => n2767);
   U2648 : AOI22_X1 port map( A1 => n5696, A2 => n6774, B1 => n2499, B2 => n566
                           , ZN => n2766);
   U2649 : NAND2_X1 port map( A1 => n2768, A2 => n2769, ZN => n2761);
   U2650 : AOI22_X1 port map( A1 => n5690, A2 => n694, B1 => n2503, B2 => n662,
                           ZN => n2769);
   U2651 : AOI22_X1 port map( A1 => n5684, A2 => n726, B1 => n2505, B2 => n598,
                           ZN => n2768);
   U2652 : NAND2_X1 port map( A1 => n2770, A2 => n2771, ZN => n2760);
   U2653 : AOI22_X1 port map( A1 => n5677, A2 => n502, B1 => n2509, B2 => n374,
                           ZN => n2771);
   U2654 : AOI22_X1 port map( A1 => n5672, A2 => n534, B1 => n2511, B2 => n342,
                           ZN => n2770);
   U2655 : NAND2_X1 port map( A1 => n2772, A2 => n2773, ZN => n3218);
   U2656 : NOR4_X1 port map( A1 => n2774, A2 => n2775, A3 => n2776, A4 => n2777
                           , ZN => n2773);
   U2657 : OAI21_X1 port map( B1 => n1434, B2 => n2460, A => n2778, ZN => n2777
                           );
   U2658 : NAND2_X1 port map( A1 => n5759, A2 => n6848, ZN => n2778);
   U2659 : OAI21_X1 port map( B1 => n6070, B2 => n2463, A => n2779, ZN => n2776
                           );
   U2660 : AOI22_X1 port map( A1 => n2465, A2 => n6696, B1 => n5750, B2 => 
                           n6976, ZN => n2779);
   U2661 : NAND2_X1 port map( A1 => n2780, A2 => n2781, ZN => n2775);
   U2662 : AOI22_X1 port map( A1 => n2469, A2 => n2819, B1 => n2470, B2 => 
                           n6916, ZN => n2781);
   U2663 : AOI22_X1 port map( A1 => n5741, A2 => n6615, B1 => n2472, B2 => 
                           n7040, ZN => n2780);
   U2665 : AOI22_X1 port map( A1 => n5735, A2 => n6731, B1 => n2478, B2 => 
                           n7008, ZN => n2785);
   U2666 : AOI22_X1 port map( A1 => n5729, A2 => n6656, B1 => n5725, B2 => 
                           n6915, ZN => n2784);
   U2667 : AOI22_X1 port map( A1 => n2481, A2 => n2230, B1 => n5720, B2 => 
                           n6763, ZN => n2783);
   U2668 : AOI22_X1 port map( A1 => n2483, A2 => n629, B1 => n5714, B2 => n469,
                           ZN => n2782);
   U2669 : NOR4_X1 port map( A1 => n2786, A2 => n2787, A3 => n2788, A4 => n2789
                           , ZN => n2772);
   U2670 : NAND2_X1 port map( A1 => n2790, A2 => n2791, ZN => n2789);
   U2671 : AOI22_X1 port map( A1 => n5711, A2 => n405, B1 => n2492, B2 => n7072
                           , ZN => n2791);
   U2672 : AOI22_X1 port map( A1 => n5705, A2 => n6807, B1 => n5935, B2 => 
                           OUT1_20_port, ZN => n2790);
   U2673 : NAND2_X1 port map( A1 => n2792, A2 => n2793, ZN => n2788);
   U2674 : AOI22_X1 port map( A1 => n5701, A2 => n437, B1 => n2497, B2 => n6950
                           , ZN => n2793);
   U2675 : AOI22_X1 port map( A1 => n5696, A2 => n6775, B1 => n2499, B2 => n565
                           , ZN => n2792);
   U2676 : NAND2_X1 port map( A1 => n2794, A2 => n2795, ZN => n2787);
   U2677 : AOI22_X1 port map( A1 => n5690, A2 => n693, B1 => n2503, B2 => n661,
                           ZN => n2795);
   U2678 : AOI22_X1 port map( A1 => n5684, A2 => n725, B1 => n2505, B2 => n597,
                           ZN => n2794);
   U2679 : NAND2_X1 port map( A1 => n2796, A2 => n2797, ZN => n2786);
   U2680 : AOI22_X1 port map( A1 => n5677, A2 => n501, B1 => n2509, B2 => n373,
                           ZN => n2797);
   U2681 : AOI22_X1 port map( A1 => n5672, A2 => n533, B1 => n2511, B2 => n341,
                           ZN => n2796);
   U2682 : NAND2_X1 port map( A1 => n2798, A2 => n2799, ZN => n3217);
   U2683 : NOR4_X1 port map( A1 => n2800, A2 => n2801, A3 => n2802, A4 => n2803
                           , ZN => n2799);
   U2684 : OAI21_X1 port map( B1 => n1435, B2 => n2460, A => n2804, ZN => n2803
                           );
   U2685 : NAND2_X1 port map( A1 => n5759, A2 => n6847, ZN => n2804);
   U2686 : OAI21_X1 port map( B1 => n6071, B2 => n2463, A => n2805, ZN => n2802
                           );
   U2687 : AOI22_X1 port map( A1 => n5753, A2 => n6695, B1 => n2466, B2 => 
                           n6975, ZN => n2805);
   U2688 : NAND2_X1 port map( A1 => n2806, A2 => n2831, ZN => n2801);
   U2689 : AOI22_X1 port map( A1 => n2469, A2 => n2818, B1 => n5744, B2 => 
                           n6914, ZN => n2831);
   U2690 : AOI22_X1 port map( A1 => n2471, A2 => n6616, B1 => n5738, B2 => 
                           n7039, ZN => n2806);
   U2692 : AOI22_X1 port map( A1 => n5735, A2 => n6730, B1 => n2478, B2 => 
                           n7007, ZN => n2835);
   U2693 : AOI22_X1 port map( A1 => n5729, A2 => n6655, B1 => n5725, B2 => 
                           n6913, ZN => n2834);
   U2694 : AOI22_X1 port map( A1 => n2481, A2 => n2225, B1 => n5720, B2 => 
                           n6762, ZN => n2833);
   U2695 : AOI22_X1 port map( A1 => n2483, A2 => n628, B1 => n5714, B2 => n468,
                           ZN => n2832);
   U2696 : NOR4_X1 port map( A1 => n2836, A2 => n2837, A3 => n2838, A4 => n2839
                           , ZN => n2798);
   U2697 : NAND2_X1 port map( A1 => n2840, A2 => n2841, ZN => n2839);
   U2698 : AOI22_X1 port map( A1 => n5711, A2 => n404, B1 => n2492, B2 => n7071
                           , ZN => n2841);
   U2699 : AOI22_X1 port map( A1 => n5705, A2 => n6808, B1 => n5935, B2 => 
                           OUT1_19_port, ZN => n2840);
   U2700 : NAND2_X1 port map( A1 => n2842, A2 => n2843, ZN => n2838);
   U2701 : AOI22_X1 port map( A1 => n5701, A2 => n436, B1 => n2497, B2 => n6951
                           , ZN => n2843);
   U2702 : AOI22_X1 port map( A1 => n5696, A2 => n6776, B1 => n2499, B2 => n564
                           , ZN => n2842);
   U2703 : NAND2_X1 port map( A1 => n2844, A2 => n2845, ZN => n2837);
   U2704 : AOI22_X1 port map( A1 => n5690, A2 => n692, B1 => n2503, B2 => n660,
                           ZN => n2845);
   U2705 : AOI22_X1 port map( A1 => n5684, A2 => n724, B1 => n2505, B2 => n596,
                           ZN => n2844);
   U2706 : NAND2_X1 port map( A1 => n2846, A2 => n2847, ZN => n2836);
   U2707 : AOI22_X1 port map( A1 => n5677, A2 => n500, B1 => n2509, B2 => n372,
                           ZN => n2847);
   U2708 : AOI22_X1 port map( A1 => n5672, A2 => n532, B1 => n2511, B2 => n340,
                           ZN => n2846);
   U2709 : NAND2_X1 port map( A1 => n2848, A2 => n2849, ZN => n3216);
   U2710 : NOR4_X1 port map( A1 => n2850, A2 => n2851, A3 => n2852, A4 => n2853
                           , ZN => n2849);
   U2711 : OAI21_X1 port map( B1 => n1436, B2 => n2460, A => n2854, ZN => n2853
                           );
   U2712 : NAND2_X1 port map( A1 => n2462, A2 => n6846, ZN => n2854);
   U2713 : OAI21_X1 port map( B1 => n6072, B2 => n2463, A => n2855, ZN => n2852
                           );
   U2714 : AOI22_X1 port map( A1 => n5753, A2 => n6694, B1 => n2466, B2 => 
                           n6974, ZN => n2855);
   U2715 : NAND2_X1 port map( A1 => n2856, A2 => n2857, ZN => n2851);
   U2716 : AOI22_X1 port map( A1 => n2469, A2 => n2817, B1 => n5744, B2 => 
                           n6912, ZN => n2857);
   U2717 : AOI22_X1 port map( A1 => n2471, A2 => n6617, B1 => n5738, B2 => 
                           n7038, ZN => n2856);
   U2719 : AOI22_X1 port map( A1 => n5735, A2 => n6729, B1 => n5732, B2 => 
                           n7006, ZN => n2861);
   U2720 : AOI22_X1 port map( A1 => n5729, A2 => n6654, B1 => n5725, B2 => 
                           n6911, ZN => n2860);
   U2721 : AOI22_X1 port map( A1 => n5723, A2 => n2220, B1 => n2482, B2 => 
                           n6761, ZN => n2859);
   U2722 : AOI22_X1 port map( A1 => n5717, A2 => n627, B1 => n2484, B2 => n467,
                           ZN => n2858);
   U2723 : NOR4_X1 port map( A1 => n2862, A2 => n2863, A3 => n2864, A4 => n2865
                           , ZN => n2848);
   U2724 : NAND2_X1 port map( A1 => n2866, A2 => n2867, ZN => n2865);
   U2725 : AOI22_X1 port map( A1 => n5711, A2 => n403, B1 => n2492, B2 => n7070
                           , ZN => n2867);
   U2726 : AOI22_X1 port map( A1 => n5705, A2 => n6809, B1 => n5935, B2 => 
                           OUT1_18_port, ZN => n2866);
   U2727 : NAND2_X1 port map( A1 => n2868, A2 => n2869, ZN => n2864);
   U2728 : AOI22_X1 port map( A1 => n5701, A2 => n435, B1 => n2497, B2 => n6952
                           , ZN => n2869);
   U2729 : AOI22_X1 port map( A1 => n5696, A2 => n6777, B1 => n2499, B2 => n563
                           , ZN => n2868);
   U2730 : NAND2_X1 port map( A1 => n2870, A2 => n2871, ZN => n2863);
   U2731 : AOI22_X1 port map( A1 => n5690, A2 => n691, B1 => n2503, B2 => n659,
                           ZN => n2871);
   U2732 : AOI22_X1 port map( A1 => n5684, A2 => n723, B1 => n2505, B2 => n595,
                           ZN => n2870);
   U2733 : NAND2_X1 port map( A1 => n2872, A2 => n2873, ZN => n2862);
   U2734 : AOI22_X1 port map( A1 => n5677, A2 => n499, B1 => n2509, B2 => n371,
                           ZN => n2873);
   U2735 : AOI22_X1 port map( A1 => n5672, A2 => n531, B1 => n2511, B2 => n339,
                           ZN => n2872);
   U2736 : NAND2_X1 port map( A1 => n2874, A2 => n2875, ZN => n3215);
   U2737 : NOR4_X1 port map( A1 => n2876, A2 => n2877, A3 => n2878, A4 => n2879
                           , ZN => n2875);
   U2738 : OAI21_X1 port map( B1 => n1437, B2 => n2460, A => n2880, ZN => n2879
                           );
   U2739 : NAND2_X1 port map( A1 => n2462, A2 => n6845, ZN => n2880);
   U2740 : OAI21_X1 port map( B1 => n5499, B2 => n2463, A => n2881, ZN => n2878
                           );
   U2741 : AOI22_X1 port map( A1 => n5753, A2 => n6693, B1 => n2466, B2 => 
                           n6973, ZN => n2881);
   U2742 : NAND2_X1 port map( A1 => n2882, A2 => n2883, ZN => n2877);
   U2743 : AOI22_X1 port map( A1 => n2469, A2 => n2816, B1 => n5744, B2 => 
                           n6910, ZN => n2883);
   U2744 : AOI22_X1 port map( A1 => n2471, A2 => n6618, B1 => n5738, B2 => 
                           n7037, ZN => n2882);
   U2746 : AOI22_X1 port map( A1 => n2477, A2 => n6728, B1 => n5732, B2 => 
                           n7005, ZN => n2887);
   U2747 : AOI22_X1 port map( A1 => n2479, A2 => n6653, B1 => n5725, B2 => 
                           n6909, ZN => n2886);
   U2748 : AOI22_X1 port map( A1 => n5723, A2 => n2215, B1 => n2482, B2 => 
                           n6760, ZN => n2885);
   U2749 : AOI22_X1 port map( A1 => n5717, A2 => n626, B1 => n2484, B2 => n466,
                           ZN => n2884);
   U2750 : NOR4_X1 port map( A1 => n2888, A2 => n2889, A3 => n2890, A4 => n2891
                           , ZN => n2874);
   U2751 : NAND2_X1 port map( A1 => n2892, A2 => n2893, ZN => n2891);
   U2752 : AOI22_X1 port map( A1 => n2491, A2 => n402, B1 => n5708, B2 => n7069
                           , ZN => n2893);
   U2753 : AOI22_X1 port map( A1 => n2493, A2 => n6810, B1 => n5935, B2 => 
                           OUT1_17_port, ZN => n2892);
   U2754 : NAND2_X1 port map( A1 => n2894, A2 => n2895, ZN => n2890);
   U2755 : AOI22_X1 port map( A1 => n5701, A2 => n434, B1 => n2497, B2 => n6953
                           , ZN => n2895);
   U2756 : AOI22_X1 port map( A1 => n2498, A2 => n6778, B1 => n5693, B2 => n562
                           , ZN => n2894);
   U2757 : NAND2_X1 port map( A1 => n2896, A2 => n2897, ZN => n2889);
   U2758 : AOI22_X1 port map( A1 => n5690, A2 => n690, B1 => n5687, B2 => n658,
                           ZN => n2897);
   U2759 : AOI22_X1 port map( A1 => n2504, A2 => n722, B1 => n5681, B2 => n594,
                           ZN => n2896);
   U2760 : NAND2_X1 port map( A1 => n2898, A2 => n2899, ZN => n2888);
   U2761 : AOI22_X1 port map( A1 => n5677, A2 => n498, B1 => n2509, B2 => n370,
                           ZN => n2899);
   U2762 : AOI22_X1 port map( A1 => n2510, A2 => n530, B1 => n5669, B2 => n338,
                           ZN => n2898);
   U2763 : NAND2_X1 port map( A1 => n2900, A2 => n2901, ZN => n3214);
   U2764 : NOR4_X1 port map( A1 => n2902, A2 => n2903, A3 => n2904, A4 => n2905
                           , ZN => n2901);
   U2765 : OAI21_X1 port map( B1 => n1438, B2 => n2460, A => n2906, ZN => n2905
                           );
   U2766 : NAND2_X1 port map( A1 => n2462, A2 => n6844, ZN => n2906);
   U2767 : OAI21_X1 port map( B1 => n6074, B2 => n2463, A => n2907, ZN => n2904
                           );
   U2768 : AOI22_X1 port map( A1 => n5753, A2 => n6692, B1 => n2466, B2 => 
                           n6972, ZN => n2907);
   U2769 : NAND2_X1 port map( A1 => n2908, A2 => n2909, ZN => n2903);
   U2770 : AOI22_X1 port map( A1 => n2469, A2 => n2815, B1 => n5744, B2 => 
                           n6908, ZN => n2909);
   U2771 : AOI22_X1 port map( A1 => n2471, A2 => n6619, B1 => n5738, B2 => 
                           n7036, ZN => n2908);
   U2773 : AOI22_X1 port map( A1 => n2477, A2 => n6727, B1 => n5732, B2 => 
                           n7004, ZN => n2913);
   U2774 : AOI22_X1 port map( A1 => n2479, A2 => n6652, B1 => n5725, B2 => 
                           n6907, ZN => n2912);
   U2775 : AOI22_X1 port map( A1 => n5723, A2 => n2210, B1 => n2482, B2 => 
                           n6759, ZN => n2911);
   U2776 : AOI22_X1 port map( A1 => n5717, A2 => n625, B1 => n2484, B2 => n465,
                           ZN => n2910);
   U2777 : NOR4_X1 port map( A1 => n2914, A2 => n2915, A3 => n2916, A4 => n2917
                           , ZN => n2900);
   U2778 : NAND2_X1 port map( A1 => n2918, A2 => n2919, ZN => n2917);
   U2779 : AOI22_X1 port map( A1 => n2491, A2 => n401, B1 => n5708, B2 => n7068
                           , ZN => n2919);
   U2780 : AOI22_X1 port map( A1 => n2493, A2 => n6811, B1 => n5935, B2 => 
                           OUT1_16_port, ZN => n2918);
   U2781 : NAND2_X1 port map( A1 => n2920, A2 => n2921, ZN => n2916);
   U2782 : AOI22_X1 port map( A1 => n5701, A2 => n433, B1 => n2497, B2 => n6954
                           , ZN => n2921);
   U2783 : AOI22_X1 port map( A1 => n2498, A2 => n6779, B1 => n5693, B2 => n561
                           , ZN => n2920);
   U2784 : NAND2_X1 port map( A1 => n2922, A2 => n2923, ZN => n2915);
   U2785 : AOI22_X1 port map( A1 => n2502, A2 => n689, B1 => n5687, B2 => n657,
                           ZN => n2923);
   U2786 : AOI22_X1 port map( A1 => n2504, A2 => n721, B1 => n5681, B2 => n593,
                           ZN => n2922);
   U2787 : NAND2_X1 port map( A1 => n2924, A2 => n2925, ZN => n2914);
   U2788 : AOI22_X1 port map( A1 => n5677, A2 => n497, B1 => n2509, B2 => n369,
                           ZN => n2925);
   U2789 : AOI22_X1 port map( A1 => n2510, A2 => n529, B1 => n5669, B2 => n337,
                           ZN => n2924);
   U2790 : NAND2_X1 port map( A1 => n2926, A2 => n2927, ZN => n3213);
   U2791 : NOR4_X1 port map( A1 => n2928, A2 => n2929, A3 => n2930, A4 => n2931
                           , ZN => n2927);
   U2792 : OAI21_X1 port map( B1 => n1439, B2 => n2460, A => n2932, ZN => n2931
                           );
   U2793 : NAND2_X1 port map( A1 => n5759, A2 => n6843, ZN => n2932);
   U2794 : OAI21_X1 port map( B1 => n6075, B2 => n2463, A => n2933, ZN => n2930
                           );
   U2795 : AOI22_X1 port map( A1 => n5753, A2 => n6691, B1 => n5750, B2 => 
                           n6971, ZN => n2933);
   U2796 : NAND2_X1 port map( A1 => n2934, A2 => n2935, ZN => n2929);
   U2797 : AOI22_X1 port map( A1 => n5745, A2 => n2814, B1 => n5744, B2 => 
                           n6906, ZN => n2935);
   U2798 : AOI22_X1 port map( A1 => n5741, A2 => n6620, B1 => n5738, B2 => 
                           n7035, ZN => n2934);
   U2800 : AOI22_X1 port map( A1 => n5735, A2 => n6726, B1 => n5732, B2 => 
                           n7003, ZN => n2939);
   U2801 : AOI22_X1 port map( A1 => n5729, A2 => n6651, B1 => n5725, B2 => 
                           n6905, ZN => n2938);
   U2802 : AOI22_X1 port map( A1 => n5723, A2 => n2205, B1 => n5720, B2 => 
                           n6758, ZN => n2937);
   U2803 : AOI22_X1 port map( A1 => n5717, A2 => n624, B1 => n5714, B2 => n464,
                           ZN => n2936);
   U2804 : NOR4_X1 port map( A1 => n2940, A2 => n2941, A3 => n2942, A4 => n2943
                           , ZN => n2926);
   U2805 : NAND2_X1 port map( A1 => n2944, A2 => n2945, ZN => n2943);
   U2806 : AOI22_X1 port map( A1 => n2491, A2 => n400, B1 => n5708, B2 => n7067
                           , ZN => n2945);
   U2807 : AOI22_X1 port map( A1 => n2493, A2 => n6812, B1 => n5935, B2 => 
                           OUT1_15_port, ZN => n2944);
   U2808 : NAND2_X1 port map( A1 => n2946, A2 => n2947, ZN => n2942);
   U2809 : AOI22_X1 port map( A1 => n5701, A2 => n432, B1 => n2497, B2 => n6955
                           , ZN => n2947);
   U2810 : AOI22_X1 port map( A1 => n2498, A2 => n6780, B1 => n5693, B2 => n560
                           , ZN => n2946);
   U2811 : NAND2_X1 port map( A1 => n2948, A2 => n2949, ZN => n2941);
   U2812 : AOI22_X1 port map( A1 => n2502, A2 => n688, B1 => n5687, B2 => n656,
                           ZN => n2949);
   U2813 : AOI22_X1 port map( A1 => n2504, A2 => n720, B1 => n5681, B2 => n592,
                           ZN => n2948);
   U2814 : NAND2_X1 port map( A1 => n2950, A2 => n2951, ZN => n2940);
   U2815 : AOI22_X1 port map( A1 => n5677, A2 => n496, B1 => n2509, B2 => n368,
                           ZN => n2951);
   U2816 : AOI22_X1 port map( A1 => n2510, A2 => n528, B1 => n5669, B2 => n336,
                           ZN => n2950);
   U2817 : NAND2_X1 port map( A1 => n2952, A2 => n2953, ZN => n3212);
   U2818 : NOR4_X1 port map( A1 => n2954, A2 => n2955, A3 => n2956, A4 => n2957
                           , ZN => n2953);
   U2819 : OAI21_X1 port map( B1 => n1440, B2 => n2460, A => n2958, ZN => n2957
                           );
   U2820 : NAND2_X1 port map( A1 => n2462, A2 => n6842, ZN => n2958);
   U2821 : OAI21_X1 port map( B1 => n6076, B2 => n2463, A => n2959, ZN => n2956
                           );
   U2822 : AOI22_X1 port map( A1 => n5753, A2 => n6690, B1 => n2466, B2 => 
                           n6904, ZN => n2959);
   U2823 : NAND2_X1 port map( A1 => n2960, A2 => n2961, ZN => n2955);
   U2824 : AOI22_X1 port map( A1 => n2469, A2 => n2813, B1 => n5744, B2 => 
                           n6903, ZN => n2961);
   U2825 : AOI22_X1 port map( A1 => n5741, A2 => n6621, B1 => n2472, B2 => 
                           n7034, ZN => n2960);
   U2827 : AOI22_X1 port map( A1 => n2477, A2 => n6725, B1 => n5732, B2 => 
                           n7002, ZN => n2965);
   U2828 : AOI22_X1 port map( A1 => n2479, A2 => n6650, B1 => n5725, B2 => 
                           n6902, ZN => n2964);
   U2829 : AOI22_X1 port map( A1 => n5723, A2 => n2200, B1 => n2482, B2 => 
                           n6757, ZN => n2963);
   U2830 : AOI22_X1 port map( A1 => n5717, A2 => n623, B1 => n2484, B2 => n463,
                           ZN => n2962);
   U2831 : NOR4_X1 port map( A1 => n2966, A2 => n2967, A3 => n2968, A4 => n2969
                           , ZN => n2952);
   U2832 : NAND2_X1 port map( A1 => n2970, A2 => n2971, ZN => n2969);
   U2833 : AOI22_X1 port map( A1 => n2491, A2 => n399, B1 => n5708, B2 => n7066
                           , ZN => n2971);
   U2834 : AOI22_X1 port map( A1 => n2493, A2 => n6813, B1 => n5935, B2 => 
                           OUT1_14_port, ZN => n2970);
   U2835 : NAND2_X1 port map( A1 => n2972, A2 => n2973, ZN => n2968);
   U2836 : AOI22_X1 port map( A1 => n5701, A2 => n431, B1 => n2497, B2 => n6956
                           , ZN => n2973);
   U2837 : AOI22_X1 port map( A1 => n2498, A2 => n6781, B1 => n5693, B2 => n559
                           , ZN => n2972);
   U2838 : NAND2_X1 port map( A1 => n2974, A2 => n2975, ZN => n2967);
   U2839 : AOI22_X1 port map( A1 => n2502, A2 => n687, B1 => n5687, B2 => n655,
                           ZN => n2975);
   U2840 : AOI22_X1 port map( A1 => n2504, A2 => n719, B1 => n5681, B2 => n591,
                           ZN => n2974);
   U2841 : NAND2_X1 port map( A1 => n2976, A2 => n2977, ZN => n2966);
   U2842 : AOI22_X1 port map( A1 => n5677, A2 => n495, B1 => n2509, B2 => n367,
                           ZN => n2977);
   U2843 : AOI22_X1 port map( A1 => n2510, A2 => n527, B1 => n5669, B2 => n335,
                           ZN => n2976);
   U2844 : NAND2_X1 port map( A1 => n2978, A2 => n2979, ZN => n3211);
   U2845 : NOR4_X1 port map( A1 => n2980, A2 => n2981, A3 => n2982, A4 => n2983
                           , ZN => n2979);
   U2846 : OAI21_X1 port map( B1 => n1441, B2 => n2460, A => n2984, ZN => n2983
                           );
   U2847 : NAND2_X1 port map( A1 => n2462, A2 => n6841, ZN => n2984);
   U2848 : OAI21_X1 port map( B1 => n6077, B2 => n2463, A => n2985, ZN => n2982
                           );
   U2849 : AOI22_X1 port map( A1 => n2465, A2 => n6689, B1 => n5750, B2 => 
                           n6901, ZN => n2985);
   U2850 : NAND2_X1 port map( A1 => n2986, A2 => n2987, ZN => n2981);
   U2851 : AOI22_X1 port map( A1 => n2469, A2 => n2812, B1 => n2470, B2 => 
                           n6900, ZN => n2987);
   U2852 : AOI22_X1 port map( A1 => n5741, A2 => n6622, B1 => n2472, B2 => 
                           n7033, ZN => n2986);
   U2854 : AOI22_X1 port map( A1 => n2477, A2 => n6724, B1 => n5732, B2 => 
                           n7001, ZN => n2991);
   U2855 : AOI22_X1 port map( A1 => n2479, A2 => n6649, B1 => n5725, B2 => 
                           n6899, ZN => n2990);
   U2856 : AOI22_X1 port map( A1 => n5723, A2 => n2195, B1 => n2482, B2 => 
                           n6756, ZN => n2989);
   U2857 : AOI22_X1 port map( A1 => n5717, A2 => n622, B1 => n2484, B2 => n462,
                           ZN => n2988);
   U2858 : NOR4_X1 port map( A1 => n2992, A2 => n2993, A3 => n2994, A4 => n2995
                           , ZN => n2978);
   U2859 : NAND2_X1 port map( A1 => n2996, A2 => n2997, ZN => n2995);
   U2860 : AOI22_X1 port map( A1 => n2491, A2 => n398, B1 => n5708, B2 => n7065
                           , ZN => n2997);
   U2861 : AOI22_X1 port map( A1 => n2493, A2 => n6814, B1 => n5935, B2 => 
                           OUT1_13_port, ZN => n2996);
   U2862 : NAND2_X1 port map( A1 => n2998, A2 => n2999, ZN => n2994);
   U2863 : AOI22_X1 port map( A1 => n5701, A2 => n430, B1 => n2497, B2 => n6957
                           , ZN => n2999);
   U2864 : AOI22_X1 port map( A1 => n2498, A2 => n6782, B1 => n5693, B2 => n558
                           , ZN => n2998);
   U2865 : NAND2_X1 port map( A1 => n3000, A2 => n3001, ZN => n2993);
   U2866 : AOI22_X1 port map( A1 => n2502, A2 => n686, B1 => n5687, B2 => n654,
                           ZN => n3001);
   U2867 : AOI22_X1 port map( A1 => n2504, A2 => n718, B1 => n5681, B2 => n590,
                           ZN => n3000);
   U2868 : NAND2_X1 port map( A1 => n3002, A2 => n3003, ZN => n2992);
   U2869 : AOI22_X1 port map( A1 => n5677, A2 => n494, B1 => n2509, B2 => n366,
                           ZN => n3003);
   U2870 : AOI22_X1 port map( A1 => n2510, A2 => n526, B1 => n5669, B2 => n334,
                           ZN => n3002);
   U2871 : NAND2_X1 port map( A1 => n3004, A2 => n3005, ZN => n3210);
   U2872 : NOR4_X1 port map( A1 => n3006, A2 => n3007, A3 => n3008, A4 => n3009
                           , ZN => n3005);
   U2873 : OAI21_X1 port map( B1 => n1442, B2 => n2460, A => n3010, ZN => n3009
                           );
   U2874 : NAND2_X1 port map( A1 => n2462, A2 => n6840, ZN => n3010);
   U2875 : OAI21_X1 port map( B1 => n6078, B2 => n2463, A => n3011, ZN => n3008
                           );
   U2876 : AOI22_X1 port map( A1 => n2465, A2 => n6688, B1 => n5750, B2 => 
                           n6898, ZN => n3011);
   U2877 : NAND2_X1 port map( A1 => n3012, A2 => n3013, ZN => n3007);
   U2878 : AOI22_X1 port map( A1 => n2469, A2 => n2811, B1 => n2470, B2 => 
                           n6897, ZN => n3013);
   U2879 : AOI22_X1 port map( A1 => n5741, A2 => n6623, B1 => n2472, B2 => 
                           n7032, ZN => n3012);
   U2881 : AOI22_X1 port map( A1 => n2477, A2 => n6723, B1 => n5732, B2 => 
                           n7000, ZN => n3017);
   U2882 : AOI22_X1 port map( A1 => n2479, A2 => n6648, B1 => n5725, B2 => 
                           n6896, ZN => n3016);
   U2883 : AOI22_X1 port map( A1 => n5723, A2 => n2190, B1 => n2482, B2 => 
                           n6755, ZN => n3015);
   U2884 : AOI22_X1 port map( A1 => n5717, A2 => n621, B1 => n2484, B2 => n461,
                           ZN => n3014);
   U2885 : NOR4_X1 port map( A1 => n3018, A2 => n3019, A3 => n3020, A4 => n3021
                           , ZN => n3004);
   U2886 : NAND2_X1 port map( A1 => n3022, A2 => n3023, ZN => n3021);
   U2887 : AOI22_X1 port map( A1 => n5711, A2 => n397, B1 => n2492, B2 => n7064
                           , ZN => n3023);
   U2888 : AOI22_X1 port map( A1 => n5705, A2 => n6815, B1 => n5934, B2 => 
                           OUT1_12_port, ZN => n3022);
   U2889 : NAND2_X1 port map( A1 => n3024, A2 => n3025, ZN => n3020);
   U2890 : AOI22_X1 port map( A1 => n5701, A2 => n429, B1 => n5697, B2 => n6958
                           , ZN => n3025);
   U2891 : AOI22_X1 port map( A1 => n5696, A2 => n6783, B1 => n5693, B2 => n557
                           , ZN => n3024);
   U2892 : NAND2_X1 port map( A1 => n3026, A2 => n3027, ZN => n3019);
   U2893 : AOI22_X1 port map( A1 => n5690, A2 => n685, B1 => n5687, B2 => n653,
                           ZN => n3027);
   U2894 : AOI22_X1 port map( A1 => n5684, A2 => n717, B1 => n5681, B2 => n589,
                           ZN => n3026);
   U2895 : NAND2_X1 port map( A1 => n3028, A2 => n3029, ZN => n3018);
   U2896 : AOI22_X1 port map( A1 => n5677, A2 => n493, B1 => n5673, B2 => n365,
                           ZN => n3029);
   U2897 : AOI22_X1 port map( A1 => n5672, A2 => n525, B1 => n5669, B2 => n333,
                           ZN => n3028);
   U2898 : NAND2_X1 port map( A1 => n3030, A2 => n3031, ZN => n3209);
   U2899 : NOR4_X1 port map( A1 => n3032, A2 => n3033, A3 => n3034, A4 => n3035
                           , ZN => n3031);
   U2900 : OAI21_X1 port map( B1 => n1443, B2 => n2460, A => n3036, ZN => n3035
                           );
   U2901 : NAND2_X1 port map( A1 => n2462, A2 => n6839, ZN => n3036);
   U2902 : OAI21_X1 port map( B1 => n6079, B2 => n2463, A => n3037, ZN => n3034
                           );
   U2903 : AOI22_X1 port map( A1 => n2465, A2 => n6687, B1 => n2466, B2 => 
                           n6895, ZN => n3037);
   U2904 : NAND2_X1 port map( A1 => n3038, A2 => n3039, ZN => n3033);
   U2905 : AOI22_X1 port map( A1 => n5745, A2 => n2810, B1 => n2470, B2 => 
                           n6894, ZN => n3039);
   U2906 : AOI22_X1 port map( A1 => n2471, A2 => n6624, B1 => n2472, B2 => 
                           n7031, ZN => n3038);
   U2908 : AOI22_X1 port map( A1 => n2477, A2 => n6722, B1 => n2478, B2 => 
                           n6999, ZN => n3043);
   U2909 : AOI22_X1 port map( A1 => n2479, A2 => n6647, B1 => n5725, B2 => 
                           n6893, ZN => n3042);
   U2910 : AOI22_X1 port map( A1 => n2481, A2 => n2185, B1 => n2482, B2 => 
                           n6754, ZN => n3041);
   U2911 : AOI22_X1 port map( A1 => n2483, A2 => n620, B1 => n2484, B2 => n460,
                           ZN => n3040);
   U2912 : NOR4_X1 port map( A1 => n3044, A2 => n3045, A3 => n3046, A4 => n3047
                           , ZN => n3030);
   U2913 : NAND2_X1 port map( A1 => n3048, A2 => n3049, ZN => n3047);
   U2914 : AOI22_X1 port map( A1 => n5711, A2 => n396, B1 => n2492, B2 => n7063
                           , ZN => n3049);
   U2915 : AOI22_X1 port map( A1 => n2493, A2 => n6816, B1 => n5934, B2 => 
                           OUT1_11_port, ZN => n3048);
   U2916 : NAND2_X1 port map( A1 => n3050, A2 => n3051, ZN => n3046);
   U2917 : AOI22_X1 port map( A1 => n5701, A2 => n428, B1 => n5697, B2 => n6959
                           , ZN => n3051);
   U2918 : AOI22_X1 port map( A1 => n2498, A2 => n6784, B1 => n2499, B2 => n556
                           , ZN => n3050);
   U2919 : NAND2_X1 port map( A1 => n3052, A2 => n3053, ZN => n3045);
   U2920 : AOI22_X1 port map( A1 => n2502, A2 => n684, B1 => n2503, B2 => n652,
                           ZN => n3053);
   U2921 : AOI22_X1 port map( A1 => n2504, A2 => n716, B1 => n2505, B2 => n588,
                           ZN => n3052);
   U2922 : NAND2_X1 port map( A1 => n3054, A2 => n3919, ZN => n3044);
   U2923 : AOI22_X1 port map( A1 => n5677, A2 => n492, B1 => n5673, B2 => n364,
                           ZN => n3919);
   U2924 : AOI22_X1 port map( A1 => n2510, A2 => n524, B1 => n2511, B2 => n332,
                           ZN => n3054);
   U2925 : NAND2_X1 port map( A1 => n3920, A2 => n3921, ZN => n3208);
   U2926 : NOR4_X1 port map( A1 => n3922, A2 => n3923, A3 => n3924, A4 => n3925
                           , ZN => n3921);
   U2927 : OAI21_X1 port map( B1 => n1444, B2 => n2460, A => n3926, ZN => n3925
                           );
   U2928 : NAND2_X1 port map( A1 => n2462, A2 => n6838, ZN => n3926);
   U2929 : OAI21_X1 port map( B1 => n6080, B2 => n2463, A => n3927, ZN => n3924
                           );
   U2930 : AOI22_X1 port map( A1 => n2465, A2 => n6686, B1 => n2466, B2 => 
                           n6892, ZN => n3927);
   U2931 : NAND2_X1 port map( A1 => n3928, A2 => n3929, ZN => n3923);
   U2932 : AOI22_X1 port map( A1 => n5745, A2 => n2809, B1 => n2470, B2 => 
                           n6891, ZN => n3929);
   U2933 : AOI22_X1 port map( A1 => n2471, A2 => n6625, B1 => n2472, B2 => 
                           n7030, ZN => n3928);
   U2935 : AOI22_X1 port map( A1 => n2477, A2 => n6721, B1 => n2478, B2 => 
                           n6998, ZN => n3933);
   U2936 : AOI22_X1 port map( A1 => n2479, A2 => n6646, B1 => n5725, B2 => 
                           n6890, ZN => n3932);
   U2937 : AOI22_X1 port map( A1 => n2481, A2 => n2180, B1 => n2482, B2 => 
                           n6753, ZN => n3931);
   U2938 : AOI22_X1 port map( A1 => n2483, A2 => n619, B1 => n2484, B2 => n459,
                           ZN => n3930);
   U2939 : NOR4_X1 port map( A1 => n3934, A2 => n3935, A3 => n3936, A4 => n3937
                           , ZN => n3920);
   U2940 : NAND2_X1 port map( A1 => n3938, A2 => n3939, ZN => n3937);
   U2941 : AOI22_X1 port map( A1 => n5711, A2 => n395, B1 => n2492, B2 => n7062
                           , ZN => n3939);
   U2942 : AOI22_X1 port map( A1 => n2493, A2 => n6817, B1 => n5934, B2 => 
                           OUT1_10_port, ZN => n3938);
   U2943 : NAND2_X1 port map( A1 => n3940, A2 => n3941, ZN => n3936);
   U2944 : AOI22_X1 port map( A1 => n5701, A2 => n427, B1 => n5697, B2 => n6960
                           , ZN => n3941);
   U2945 : AOI22_X1 port map( A1 => n2498, A2 => n6785, B1 => n2499, B2 => n555
                           , ZN => n3940);
   U2946 : NAND2_X1 port map( A1 => n3942, A2 => n3943, ZN => n3935);
   U2947 : AOI22_X1 port map( A1 => n2502, A2 => n683, B1 => n2503, B2 => n651,
                           ZN => n3943);
   U2948 : AOI22_X1 port map( A1 => n2504, A2 => n715, B1 => n2505, B2 => n587,
                           ZN => n3942);
   U2949 : NAND2_X1 port map( A1 => n3944, A2 => n3945, ZN => n3934);
   U2950 : AOI22_X1 port map( A1 => n5677, A2 => n491, B1 => n5673, B2 => n363,
                           ZN => n3945);
   U2951 : AOI22_X1 port map( A1 => n2510, A2 => n523, B1 => n2511, B2 => n331,
                           ZN => n3944);
   U2952 : NAND2_X1 port map( A1 => n3946, A2 => n3947, ZN => n3207);
   U2953 : NOR4_X1 port map( A1 => n3948, A2 => n3949, A3 => n3950, A4 => n3951
                           , ZN => n3947);
   U2954 : OAI21_X1 port map( B1 => n1445, B2 => n2460, A => n3952, ZN => n3951
                           );
   U2955 : NAND2_X1 port map( A1 => n2462, A2 => n6837, ZN => n3952);
   U2956 : OAI21_X1 port map( B1 => n5523, B2 => n2463, A => n3953, ZN => n3950
                           );
   U2957 : AOI22_X1 port map( A1 => n2465, A2 => n6685, B1 => n2466, B2 => 
                           n6889, ZN => n3953);
   U2958 : NAND2_X1 port map( A1 => n3954, A2 => n3955, ZN => n3949);
   U2959 : AOI22_X1 port map( A1 => n5745, A2 => n2808, B1 => n2470, B2 => 
                           n6888, ZN => n3955);
   U2960 : AOI22_X1 port map( A1 => n2471, A2 => n6626, B1 => n2472, B2 => 
                           n7029, ZN => n3954);
   U2962 : AOI22_X1 port map( A1 => n2477, A2 => n6720, B1 => n2478, B2 => 
                           n6997, ZN => n3959);
   U2963 : AOI22_X1 port map( A1 => n2479, A2 => n6645, B1 => n5725, B2 => 
                           n6887, ZN => n3958);
   U2964 : AOI22_X1 port map( A1 => n2481, A2 => n2175, B1 => n2482, B2 => 
                           n6752, ZN => n3957);
   U2965 : AOI22_X1 port map( A1 => n2483, A2 => n618, B1 => n2484, B2 => n458,
                           ZN => n3956);
   U2966 : NOR4_X1 port map( A1 => n3960, A2 => n3961, A3 => n3962, A4 => n3963
                           , ZN => n3946);
   U2967 : NAND2_X1 port map( A1 => n3964, A2 => n3965, ZN => n3963);
   U2968 : AOI22_X1 port map( A1 => n5711, A2 => n394, B1 => n2492, B2 => n7061
                           , ZN => n3965);
   U2969 : AOI22_X1 port map( A1 => n2493, A2 => n6818, B1 => n5934, B2 => 
                           OUT1_9_port, ZN => n3964);
   U2970 : NAND2_X1 port map( A1 => n3966, A2 => n3967, ZN => n3962);
   U2971 : AOI22_X1 port map( A1 => n5701, A2 => n426, B1 => n5697, B2 => n6961
                           , ZN => n3967);
   U2972 : AOI22_X1 port map( A1 => n2498, A2 => n6786, B1 => n2499, B2 => n554
                           , ZN => n3966);
   U2973 : NAND2_X1 port map( A1 => n3968, A2 => n3969, ZN => n3961);
   U2974 : AOI22_X1 port map( A1 => n2502, A2 => n682, B1 => n2503, B2 => n650,
                           ZN => n3969);
   U2975 : AOI22_X1 port map( A1 => n2504, A2 => n714, B1 => n2505, B2 => n586,
                           ZN => n3968);
   U2976 : NAND2_X1 port map( A1 => n3970, A2 => n3971, ZN => n3960);
   U2977 : AOI22_X1 port map( A1 => n5677, A2 => n490, B1 => n5673, B2 => n362,
                           ZN => n3971);
   U2978 : AOI22_X1 port map( A1 => n2510, A2 => n522, B1 => n2511, B2 => n330,
                           ZN => n3970);
   U2979 : NAND2_X1 port map( A1 => n3972, A2 => n3973, ZN => n3206);
   U2980 : NOR4_X1 port map( A1 => n3974, A2 => n3975, A3 => n3976, A4 => n3977
                           , ZN => n3973);
   U2981 : OAI21_X1 port map( B1 => n1446, B2 => n2460, A => n3978, ZN => n3977
                           );
   U2982 : NAND2_X1 port map( A1 => n2462, A2 => n6836, ZN => n3978);
   U2983 : OAI21_X1 port map( B1 => n6082, B2 => n2463, A => n3979, ZN => n3976
                           );
   U2984 : AOI22_X1 port map( A1 => n2465, A2 => n6684, B1 => n2466, B2 => 
                           n6886, ZN => n3979);
   U2985 : NAND2_X1 port map( A1 => n3980, A2 => n3981, ZN => n3975);
   U2986 : AOI22_X1 port map( A1 => n5745, A2 => n2807, B1 => n2470, B2 => 
                           n6885, ZN => n3981);
   U2987 : AOI22_X1 port map( A1 => n2471, A2 => n6627, B1 => n2472, B2 => 
                           n7028, ZN => n3980);
   U2989 : AOI22_X1 port map( A1 => n2477, A2 => n6719, B1 => n2478, B2 => 
                           n6996, ZN => n3985);
   U2990 : AOI22_X1 port map( A1 => n2479, A2 => n6644, B1 => n5725, B2 => 
                           n6884, ZN => n3984);
   U2991 : AOI22_X1 port map( A1 => n2481, A2 => n2170, B1 => n2482, B2 => 
                           n6751, ZN => n3983);
   U2992 : AOI22_X1 port map( A1 => n2483, A2 => n617, B1 => n2484, B2 => n457,
                           ZN => n3982);
   U2993 : NOR4_X1 port map( A1 => n3986, A2 => n3987, A3 => n3988, A4 => n3989
                           , ZN => n3972);
   U2994 : NAND2_X1 port map( A1 => n3990, A2 => n3991, ZN => n3989);
   U2995 : AOI22_X1 port map( A1 => n5711, A2 => n393, B1 => n2492, B2 => n7060
                           , ZN => n3991);
   U2996 : AOI22_X1 port map( A1 => n2493, A2 => n6819, B1 => n5934, B2 => 
                           OUT1_8_port, ZN => n3990);
   U2997 : NAND2_X1 port map( A1 => n3992, A2 => n3993, ZN => n3988);
   U2998 : AOI22_X1 port map( A1 => n5701, A2 => n425, B1 => n5697, B2 => n6962
                           , ZN => n3993);
   U2999 : AOI22_X1 port map( A1 => n2498, A2 => n6787, B1 => n2499, B2 => n553
                           , ZN => n3992);
   U3000 : NAND2_X1 port map( A1 => n3994, A2 => n3995, ZN => n3987);
   U3001 : AOI22_X1 port map( A1 => n2502, A2 => n681, B1 => n2503, B2 => n649,
                           ZN => n3995);
   U3002 : AOI22_X1 port map( A1 => n2504, A2 => n713, B1 => n2505, B2 => n585,
                           ZN => n3994);
   U3003 : NAND2_X1 port map( A1 => n3996, A2 => n3997, ZN => n3986);
   U3004 : AOI22_X1 port map( A1 => n5677, A2 => n489, B1 => n5673, B2 => n361,
                           ZN => n3997);
   U3005 : AOI22_X1 port map( A1 => n2510, A2 => n521, B1 => n2511, B2 => n329,
                           ZN => n3996);
   U3006 : NAND2_X1 port map( A1 => n4190, A2 => n4191, ZN => n3205);
   U3007 : NOR4_X1 port map( A1 => n4192, A2 => n4193, A3 => n4194, A4 => n4195
                           , ZN => n4191);
   U3008 : OAI21_X1 port map( B1 => n1447, B2 => n2460, A => n4196, ZN => n4195
                           );
   U3009 : NAND2_X1 port map( A1 => n2462, A2 => n6835, ZN => n4196);
   U3010 : OAI21_X1 port map( B1 => n6083, B2 => n2463, A => n4197, ZN => n4194
                           );
   U3011 : AOI22_X1 port map( A1 => n2465, A2 => n6683, B1 => n2466, B2 => 
                           n6883, ZN => n4197);
   U3012 : NAND2_X1 port map( A1 => n4198, A2 => n4199, ZN => n4193);
   U3013 : AOI22_X1 port map( A1 => n5745, A2 => n6675, B1 => n2470, B2 => 
                           n6882, ZN => n4199);
   U3014 : AOI22_X1 port map( A1 => n2471, A2 => n6628, B1 => n2472, B2 => 
                           n7027, ZN => n4198);
   U3016 : AOI22_X1 port map( A1 => n2477, A2 => n6718, B1 => n2478, B2 => 
                           n6995, ZN => n4203);
   U3017 : AOI22_X1 port map( A1 => n2479, A2 => n6643, B1 => n5725, B2 => 
                           n6881, ZN => n4202);
   U3018 : AOI22_X1 port map( A1 => n2481, A2 => n2165, B1 => n2482, B2 => 
                           n6750, ZN => n4201);
   U3019 : AOI22_X1 port map( A1 => n2483, A2 => n616, B1 => n2484, B2 => n456,
                           ZN => n4200);
   U3020 : NOR4_X1 port map( A1 => n4204, A2 => n4205, A3 => n4206, A4 => n4207
                           , ZN => n4190);
   U3021 : NAND2_X1 port map( A1 => n4208, A2 => n4209, ZN => n4207);
   U3022 : AOI22_X1 port map( A1 => n5711, A2 => n392, B1 => n2492, B2 => n7059
                           , ZN => n4209);
   U3023 : AOI22_X1 port map( A1 => n2493, A2 => n6820, B1 => n5934, B2 => 
                           OUT1_7_port, ZN => n4208);
   U3024 : NAND2_X1 port map( A1 => n4210, A2 => n4211, ZN => n4206);
   U3025 : AOI22_X1 port map( A1 => n5701, A2 => n424, B1 => n5697, B2 => n6963
                           , ZN => n4211);
   U3026 : AOI22_X1 port map( A1 => n2498, A2 => n6788, B1 => n2499, B2 => n552
                           , ZN => n4210);
   U3027 : NAND2_X1 port map( A1 => n4212, A2 => n4213, ZN => n4205);
   U3028 : AOI22_X1 port map( A1 => n2502, A2 => n680, B1 => n2503, B2 => n648,
                           ZN => n4213);
   U3029 : AOI22_X1 port map( A1 => n2504, A2 => n712, B1 => n2505, B2 => n584,
                           ZN => n4212);
   U3030 : NAND2_X1 port map( A1 => n4214, A2 => n4215, ZN => n4204);
   U3031 : AOI22_X1 port map( A1 => n5677, A2 => n488, B1 => n5673, B2 => n360,
                           ZN => n4215);
   U3032 : AOI22_X1 port map( A1 => n2510, A2 => n520, B1 => n2511, B2 => n328,
                           ZN => n4214);
   U3033 : NAND2_X1 port map( A1 => n4216, A2 => n4217, ZN => n3204);
   U3034 : NOR4_X1 port map( A1 => n4218, A2 => n4219, A3 => n4220, A4 => n4221
                           , ZN => n4217);
   U3035 : OAI21_X1 port map( B1 => n1448, B2 => n2460, A => n4222, ZN => n4221
                           );
   U3036 : NAND2_X1 port map( A1 => n2462, A2 => n6834, ZN => n4222);
   U3037 : OAI21_X1 port map( B1 => n6084, B2 => n2463, A => n4223, ZN => n4220
                           );
   U3038 : AOI22_X1 port map( A1 => n2465, A2 => n6682, B1 => n2466, B2 => 
                           n6880, ZN => n4223);
   U3039 : NAND2_X1 port map( A1 => n4224, A2 => n4225, ZN => n4219);
   U3040 : AOI22_X1 port map( A1 => n5745, A2 => n6674, B1 => n2470, B2 => 
                           n6879, ZN => n4225);
   U3041 : AOI22_X1 port map( A1 => n2471, A2 => n6629, B1 => n2472, B2 => 
                           n7026, ZN => n4224);
   U3043 : AOI22_X1 port map( A1 => n2477, A2 => n6717, B1 => n2478, B2 => 
                           n6994, ZN => n4229);
   U3044 : AOI22_X1 port map( A1 => n2479, A2 => n6642, B1 => n5725, B2 => 
                           n6878, ZN => n4228);
   U3045 : AOI22_X1 port map( A1 => n2481, A2 => n2160, B1 => n2482, B2 => 
                           n6749, ZN => n4227);
   U3046 : AOI22_X1 port map( A1 => n2483, A2 => n615, B1 => n2484, B2 => n455,
                           ZN => n4226);
   U3047 : NOR4_X1 port map( A1 => n4230, A2 => n4231, A3 => n4232, A4 => n4233
                           , ZN => n4216);
   U3048 : NAND2_X1 port map( A1 => n4234, A2 => n4235, ZN => n4233);
   U3049 : AOI22_X1 port map( A1 => n5711, A2 => n391, B1 => n2492, B2 => n7058
                           , ZN => n4235);
   U3050 : AOI22_X1 port map( A1 => n2493, A2 => n6821, B1 => n5934, B2 => 
                           OUT1_6_port, ZN => n4234);
   U3051 : NAND2_X1 port map( A1 => n4236, A2 => n4237, ZN => n4232);
   U3052 : AOI22_X1 port map( A1 => n5701, A2 => n423, B1 => n5697, B2 => n6964
                           , ZN => n4237);
   U3053 : AOI22_X1 port map( A1 => n2498, A2 => n6789, B1 => n2499, B2 => n551
                           , ZN => n4236);
   U3054 : NAND2_X1 port map( A1 => n4238, A2 => n4239, ZN => n4231);
   U3055 : AOI22_X1 port map( A1 => n2502, A2 => n679, B1 => n2503, B2 => n647,
                           ZN => n4239);
   U3056 : AOI22_X1 port map( A1 => n2504, A2 => n711, B1 => n2505, B2 => n583,
                           ZN => n4238);
   U3057 : NAND2_X1 port map( A1 => n4240, A2 => n4241, ZN => n4230);
   U3058 : AOI22_X1 port map( A1 => n5677, A2 => n487, B1 => n5673, B2 => n359,
                           ZN => n4241);
   U3059 : AOI22_X1 port map( A1 => n2510, A2 => n519, B1 => n2511, B2 => n327,
                           ZN => n4240);
   U3060 : NAND2_X1 port map( A1 => n4242, A2 => n4243, ZN => n3203);
   U3061 : NOR4_X1 port map( A1 => n4244, A2 => n4245, A3 => n4246, A4 => n4247
                           , ZN => n4243);
   U3062 : OAI21_X1 port map( B1 => n1449, B2 => n2460, A => n4248, ZN => n4247
                           );
   U3063 : NAND2_X1 port map( A1 => n5759, A2 => n6833, ZN => n4248);
   U3064 : OAI21_X1 port map( B1 => n6085, B2 => n2463, A => n4249, ZN => n4246
                           );
   U3065 : AOI22_X1 port map( A1 => n5753, A2 => n6681, B1 => n5750, B2 => 
                           n6877, ZN => n4249);
   U3066 : NAND2_X1 port map( A1 => n4250, A2 => n4251, ZN => n4245);
   U3067 : AOI22_X1 port map( A1 => n5745, A2 => n6673, B1 => n2470, B2 => 
                           n6876, ZN => n4251);
   U3068 : AOI22_X1 port map( A1 => n5741, A2 => n6630, B1 => n5738, B2 => 
                           n7025, ZN => n4250);
   U3070 : AOI22_X1 port map( A1 => n5735, A2 => n6716, B1 => n2478, B2 => 
                           n6993, ZN => n4255);
   U3071 : AOI22_X1 port map( A1 => n5729, A2 => n6641, B1 => n2480, B2 => 
                           n6875, ZN => n4254);
   U3072 : AOI22_X1 port map( A1 => n5723, A2 => n2155, B1 => n5720, B2 => 
                           n6748, ZN => n4253);
   U3073 : AOI22_X1 port map( A1 => n5717, A2 => n614, B1 => n5714, B2 => n454,
                           ZN => n4252);
   U3074 : NOR4_X1 port map( A1 => n4256, A2 => n4257, A3 => n4258, A4 => n4259
                           , ZN => n4242);
   U3075 : NAND2_X1 port map( A1 => n4260, A2 => n4261, ZN => n4259);
   U3076 : AOI22_X1 port map( A1 => n2491, A2 => n390, B1 => n5708, B2 => n7057
                           , ZN => n4261);
   U3077 : AOI22_X1 port map( A1 => n5705, A2 => n6822, B1 => n5934, B2 => 
                           OUT1_5_port, ZN => n4260);
   U3078 : NAND2_X1 port map( A1 => n4262, A2 => n4263, ZN => n4258);
   U3079 : AOI22_X1 port map( A1 => n5701, A2 => n422, B1 => n5697, B2 => n6965
                           , ZN => n4263);
   U3080 : AOI22_X1 port map( A1 => n5696, A2 => n6790, B1 => n5693, B2 => n550
                           , ZN => n4262);
   U3081 : NAND2_X1 port map( A1 => n4264, A2 => n4265, ZN => n4257);
   U3082 : AOI22_X1 port map( A1 => n2502, A2 => n678, B1 => n5687, B2 => n646,
                           ZN => n4265);
   U3083 : AOI22_X1 port map( A1 => n5684, A2 => n710, B1 => n5681, B2 => n582,
                           ZN => n4264);
   U3084 : NAND2_X1 port map( A1 => n4266, A2 => n4267, ZN => n4256);
   U3085 : AOI22_X1 port map( A1 => n5677, A2 => n486, B1 => n5673, B2 => n358,
                           ZN => n4267);
   U3086 : AOI22_X1 port map( A1 => n5672, A2 => n518, B1 => n5669, B2 => n326,
                           ZN => n4266);
   U3087 : NAND2_X1 port map( A1 => n4268, A2 => n4269, ZN => n3202);
   U3088 : NOR4_X1 port map( A1 => n4270, A2 => n4271, A3 => n4272, A4 => n4273
                           , ZN => n4269);
   U3089 : OAI21_X1 port map( B1 => n1450, B2 => n2460, A => n4274, ZN => n4273
                           );
   U3090 : NAND2_X1 port map( A1 => n5759, A2 => n6832, ZN => n4274);
   U3091 : OAI21_X1 port map( B1 => n6086, B2 => n2463, A => n4275, ZN => n4272
                           );
   U3092 : AOI22_X1 port map( A1 => n5753, A2 => n6680, B1 => n5750, B2 => 
                           n6874, ZN => n4275);
   U3093 : NAND2_X1 port map( A1 => n4276, A2 => n4277, ZN => n4271);
   U3094 : AOI22_X1 port map( A1 => n5745, A2 => n6672, B1 => n5744, B2 => 
                           n6873, ZN => n4277);
   U3095 : AOI22_X1 port map( A1 => n5741, A2 => n6631, B1 => n5738, B2 => 
                           n7024, ZN => n4276);
   U3097 : AOI22_X1 port map( A1 => n5735, A2 => n6715, B1 => n5732, B2 => 
                           n6992, ZN => n4281);
   U3098 : AOI22_X1 port map( A1 => n5729, A2 => n6640, B1 => n2480, B2 => 
                           n6872, ZN => n4280);
   U3099 : AOI22_X1 port map( A1 => n5723, A2 => n2150, B1 => n5720, B2 => 
                           n6747, ZN => n4279);
   U3100 : AOI22_X1 port map( A1 => n5717, A2 => n613, B1 => n5714, B2 => n453,
                           ZN => n4278);
   U3101 : NOR4_X1 port map( A1 => n4282, A2 => n4283, A3 => n4284, A4 => n4285
                           , ZN => n4268);
   U3102 : NAND2_X1 port map( A1 => n4286, A2 => n4287, ZN => n4285);
   U3103 : AOI22_X1 port map( A1 => n2491, A2 => n389, B1 => n5708, B2 => n7056
                           , ZN => n4287);
   U3104 : AOI22_X1 port map( A1 => n5705, A2 => n6823, B1 => n5934, B2 => 
                           OUT1_4_port, ZN => n4286);
   U3105 : NAND2_X1 port map( A1 => n4288, A2 => n4289, ZN => n4284);
   U3106 : AOI22_X1 port map( A1 => n2496, A2 => n421, B1 => n5697, B2 => n6966
                           , ZN => n4289);
   U3107 : AOI22_X1 port map( A1 => n5696, A2 => n6791, B1 => n5693, B2 => n549
                           , ZN => n4288);
   U3108 : NAND2_X1 port map( A1 => n4290, A2 => n4291, ZN => n4283);
   U3109 : AOI22_X1 port map( A1 => n5690, A2 => n677, B1 => n5687, B2 => n645,
                           ZN => n4291);
   U3110 : AOI22_X1 port map( A1 => n5684, A2 => n709, B1 => n5681, B2 => n581,
                           ZN => n4290);
   U3111 : NAND2_X1 port map( A1 => n4292, A2 => n4293, ZN => n4282);
   U3112 : AOI22_X1 port map( A1 => n2508, A2 => n485, B1 => n5673, B2 => n357,
                           ZN => n4293);
   U3113 : AOI22_X1 port map( A1 => n5672, A2 => n517, B1 => n5669, B2 => n325,
                           ZN => n4292);
   U3114 : NAND2_X1 port map( A1 => n4294, A2 => n4295, ZN => n3201);
   U3115 : NOR4_X1 port map( A1 => n4296, A2 => n4297, A3 => n4298, A4 => n4299
                           , ZN => n4295);
   U3116 : OAI21_X1 port map( B1 => n1451, B2 => n5762, A => n4300, ZN => n4299
                           );
   U3117 : NAND2_X1 port map( A1 => n5759, A2 => n6831, ZN => n4300);
   U3118 : OAI21_X1 port map( B1 => n6087, B2 => n5756, A => n4301, ZN => n4298
                           );
   U3119 : AOI22_X1 port map( A1 => n5753, A2 => n6679, B1 => n5750, B2 => 
                           n6871, ZN => n4301);
   U3120 : NAND2_X1 port map( A1 => n4302, A2 => n4303, ZN => n4297);
   U3121 : AOI22_X1 port map( A1 => n5745, A2 => n6671, B1 => n5744, B2 => 
                           n6870, ZN => n4303);
   U3122 : AOI22_X1 port map( A1 => n5741, A2 => n6632, B1 => n5738, B2 => 
                           n7023, ZN => n4302);
   U3124 : AOI22_X1 port map( A1 => n5735, A2 => n6714, B1 => n5732, B2 => 
                           n6991, ZN => n4307);
   U3125 : AOI22_X1 port map( A1 => n5729, A2 => n6639, B1 => n2480, B2 => 
                           n6869, ZN => n4306);
   U3126 : AOI22_X1 port map( A1 => n5723, A2 => n2145, B1 => n5720, B2 => 
                           n6746, ZN => n4305);
   U3127 : AOI22_X1 port map( A1 => n5717, A2 => n612, B1 => n5714, B2 => n452,
                           ZN => n4304);
   U3128 : NOR4_X1 port map( A1 => n4308, A2 => n4309, A3 => n4310, A4 => n4311
                           , ZN => n4294);
   U3129 : NAND2_X1 port map( A1 => n4312, A2 => n4313, ZN => n4311);
   U3130 : AOI22_X1 port map( A1 => n2491, A2 => n388, B1 => n5708, B2 => n7055
                           , ZN => n4313);
   U3131 : AOI22_X1 port map( A1 => n5705, A2 => n6824, B1 => n5934, B2 => 
                           OUT1_3_port, ZN => n4312);
   U3132 : NAND2_X1 port map( A1 => n4314, A2 => n4315, ZN => n4310);
   U3133 : AOI22_X1 port map( A1 => n2496, A2 => n420, B1 => n5697, B2 => n6967
                           , ZN => n4315);
   U3134 : AOI22_X1 port map( A1 => n5696, A2 => n6792, B1 => n5693, B2 => n548
                           , ZN => n4314);
   U3135 : NAND2_X1 port map( A1 => n4316, A2 => n4317, ZN => n4309);
   U3136 : AOI22_X1 port map( A1 => n5690, A2 => n676, B1 => n5687, B2 => n644,
                           ZN => n4317);
   U3137 : AOI22_X1 port map( A1 => n5684, A2 => n708, B1 => n5681, B2 => n580,
                           ZN => n4316);
   U3138 : NAND2_X1 port map( A1 => n4318, A2 => n4319, ZN => n4308);
   U3139 : AOI22_X1 port map( A1 => n2508, A2 => n484, B1 => n5673, B2 => n356,
                           ZN => n4319);
   U3140 : AOI22_X1 port map( A1 => n5672, A2 => n516, B1 => n5669, B2 => n324,
                           ZN => n4318);
   U3141 : NAND2_X1 port map( A1 => n4320, A2 => n4321, ZN => n3200);
   U3142 : NOR4_X1 port map( A1 => n4322, A2 => n4323, A3 => n4324, A4 => n4325
                           , ZN => n4321);
   U3143 : OAI21_X1 port map( B1 => n1452, B2 => n5762, A => n4326, ZN => n4325
                           );
   U3144 : NAND2_X1 port map( A1 => n5759, A2 => n6830, ZN => n4326);
   U3145 : OAI21_X1 port map( B1 => n6088, B2 => n5756, A => n4327, ZN => n4324
                           );
   U3146 : AOI22_X1 port map( A1 => n5753, A2 => n6678, B1 => n5750, B2 => 
                           n6868, ZN => n4327);
   U3147 : NAND2_X1 port map( A1 => n4328, A2 => n4329, ZN => n4323);
   U3148 : AOI22_X1 port map( A1 => n5745, A2 => n6670, B1 => n5744, B2 => 
                           n6867, ZN => n4329);
   U3149 : AOI22_X1 port map( A1 => n5741, A2 => n6633, B1 => n5738, B2 => 
                           n7022, ZN => n4328);
   U3151 : AOI22_X1 port map( A1 => n5735, A2 => n6713, B1 => n5732, B2 => 
                           n6990, ZN => n4333);
   U3152 : AOI22_X1 port map( A1 => n5729, A2 => n6638, B1 => n2480, B2 => 
                           n6866, ZN => n4332);
   U3153 : AOI22_X1 port map( A1 => n5723, A2 => n2140, B1 => n5720, B2 => 
                           n6745, ZN => n4331);
   U3154 : AOI22_X1 port map( A1 => n5717, A2 => n611, B1 => n5714, B2 => n451,
                           ZN => n4330);
   U3155 : NOR4_X1 port map( A1 => n4334, A2 => n4335, A3 => n4336, A4 => n4337
                           , ZN => n4320);
   U3156 : NAND2_X1 port map( A1 => n4338, A2 => n4339, ZN => n4337);
   U3157 : AOI22_X1 port map( A1 => n2491, A2 => n387, B1 => n5708, B2 => n7054
                           , ZN => n4339);
   U3158 : AOI22_X1 port map( A1 => n5705, A2 => n6825, B1 => n5934, B2 => 
                           OUT1_2_port, ZN => n4338);
   U3159 : NAND2_X1 port map( A1 => n4340, A2 => n4341, ZN => n4336);
   U3160 : AOI22_X1 port map( A1 => n2496, A2 => n419, B1 => n5697, B2 => n6968
                           , ZN => n4341);
   U3161 : AOI22_X1 port map( A1 => n5696, A2 => n6793, B1 => n5693, B2 => n547
                           , ZN => n4340);
   U3162 : NAND2_X1 port map( A1 => n4342, A2 => n4343, ZN => n4335);
   U3163 : AOI22_X1 port map( A1 => n5690, A2 => n675, B1 => n5687, B2 => n643,
                           ZN => n4343);
   U3164 : AOI22_X1 port map( A1 => n5684, A2 => n707, B1 => n5681, B2 => n579,
                           ZN => n4342);
   U3165 : NAND2_X1 port map( A1 => n4344, A2 => n4345, ZN => n4334);
   U3166 : AOI22_X1 port map( A1 => n2508, A2 => n483, B1 => n5673, B2 => n355,
                           ZN => n4345);
   U3167 : AOI22_X1 port map( A1 => n5672, A2 => n515, B1 => n5669, B2 => n323,
                           ZN => n4344);
   U3168 : NAND2_X1 port map( A1 => n4346, A2 => n4347, ZN => n3199);
   U3169 : NOR4_X1 port map( A1 => n4348, A2 => n4349, A3 => n4350, A4 => n4351
                           , ZN => n4347);
   U3170 : OAI21_X1 port map( B1 => n1453, B2 => n5762, A => n4352, ZN => n4351
                           );
   U3171 : NAND2_X1 port map( A1 => n5759, A2 => n6829, ZN => n4352);
   U3172 : OAI21_X1 port map( B1 => n6089, B2 => n5756, A => n4353, ZN => n4350
                           );
   U3173 : AOI22_X1 port map( A1 => n5753, A2 => n6677, B1 => n5750, B2 => 
                           n6865, ZN => n4353);
   U3174 : NAND2_X1 port map( A1 => n4354, A2 => n4355, ZN => n4349);
   U3175 : AOI22_X1 port map( A1 => n5745, A2 => n6669, B1 => n5744, B2 => 
                           n6864, ZN => n4355);
   U3176 : AOI22_X1 port map( A1 => n5741, A2 => n6634, B1 => n5738, B2 => 
                           n7021, ZN => n4354);
   U3178 : AOI22_X1 port map( A1 => n5735, A2 => n6712, B1 => n5732, B2 => 
                           n6989, ZN => n4359);
   U3179 : AOI22_X1 port map( A1 => n5729, A2 => n6637, B1 => n2480, B2 => 
                           n6863, ZN => n4358);
   U3180 : AOI22_X1 port map( A1 => n5723, A2 => n2135, B1 => n5720, B2 => 
                           n6744, ZN => n4357);
   U3181 : AOI22_X1 port map( A1 => n5717, A2 => n610, B1 => n5714, B2 => n450,
                           ZN => n4356);
   U3182 : NOR4_X1 port map( A1 => n4360, A2 => n4361, A3 => n4362, A4 => n4363
                           , ZN => n4346);
   U3183 : NAND2_X1 port map( A1 => n4364, A2 => n4365, ZN => n4363);
   U3184 : AOI22_X1 port map( A1 => n2491, A2 => n386, B1 => n5708, B2 => n7053
                           , ZN => n4365);
   U3185 : AOI22_X1 port map( A1 => n5705, A2 => n6826, B1 => n5934, B2 => 
                           OUT1_1_port, ZN => n4364);
   U3186 : NAND2_X1 port map( A1 => n4366, A2 => n4367, ZN => n4362);
   U3187 : AOI22_X1 port map( A1 => n2496, A2 => n418, B1 => n5697, B2 => n6969
                           , ZN => n4367);
   U3188 : AOI22_X1 port map( A1 => n5696, A2 => n6794, B1 => n5693, B2 => n546
                           , ZN => n4366);
   U3189 : NAND2_X1 port map( A1 => n4368, A2 => n4369, ZN => n4361);
   U3190 : AOI22_X1 port map( A1 => n5690, A2 => n674, B1 => n5687, B2 => n642,
                           ZN => n4369);
   U3191 : AOI22_X1 port map( A1 => n5684, A2 => n706, B1 => n5681, B2 => n578,
                           ZN => n4368);
   U3192 : NAND2_X1 port map( A1 => n4370, A2 => n4371, ZN => n4360);
   U3193 : AOI22_X1 port map( A1 => n2508, A2 => n482, B1 => n5673, B2 => n354,
                           ZN => n4371);
   U3194 : AOI22_X1 port map( A1 => n5672, A2 => n514, B1 => n5669, B2 => n322,
                           ZN => n4370);
   U3195 : NAND2_X1 port map( A1 => n4372, A2 => n4373, ZN => n3198);
   U3196 : NOR4_X1 port map( A1 => n4374, A2 => n4375, A3 => n4376, A4 => n4377
                           , ZN => n4373);
   U3197 : OAI21_X1 port map( B1 => n1454, B2 => n5762, A => n4378, ZN => n4377
                           );
   U3198 : NAND2_X1 port map( A1 => n5759, A2 => n6828, ZN => n4378);
   U3199 : NOR2_X1 port map( A1 => n4379, A2 => n4380, ZN => n2462);
   U3200 : OR2_X1 port map( A1 => n4379, A2 => n4381, ZN => n2460);
   U3201 : OAI21_X1 port map( B1 => n6090, B2 => n5756, A => n4382, ZN => n4376
                           );
   U3202 : AOI22_X1 port map( A1 => n5753, A2 => n6676, B1 => n5750, B2 => 
                           n6862, ZN => n4382);
   U3203 : NOR2_X1 port map( A1 => n4381, A2 => n4383, ZN => n2466);
   U3204 : NOR2_X1 port map( A1 => n4383, A2 => n4380, ZN => n2465);
   U3205 : NAND2_X1 port map( A1 => n4384, A2 => n4385, ZN => n2463);
   U3206 : NOR4_X1 port map( A1 => n6603, A2 => n4386, A3 => n4387, A4 => n4388
                           , ZN => n4385);
   U3207 : NOR3_X1 port map( A1 => n4389, A2 => n4390, A3 => n4391, ZN => n4384
                           );
   U3208 : NAND2_X1 port map( A1 => n4392, A2 => n4393, ZN => n4375);
   U3209 : AOI22_X1 port map( A1 => n5745, A2 => n6668, B1 => n5744, B2 => 
                           n6861, ZN => n4393);
   U3210 : NOR2_X1 port map( A1 => n4394, A2 => n4395, ZN => n2470);
   U3211 : NOR2_X1 port map( A1 => n4395, A2 => n4396, ZN => n2469);
   U3212 : AOI22_X1 port map( A1 => n5741, A2 => n6635, B1 => n5738, B2 => 
                           n7020, ZN => n4392);
   U3213 : NOR2_X1 port map( A1 => n4397, A2 => n4383, ZN => n2472);
   U3214 : NOR2_X1 port map( A1 => n4395, A2 => n4381, ZN => n2471);
   U3216 : AOI22_X1 port map( A1 => n5735, A2 => n6711, B1 => n5732, B2 => 
                           n6988, ZN => n4401);
   U3217 : NOR2_X1 port map( A1 => n4402, A2 => n4379, ZN => n2478);
   U3218 : NOR2_X1 port map( A1 => n4403, A2 => n4394, ZN => n2477);
   U3219 : AOI22_X1 port map( A1 => n5729, A2 => n6636, B1 => n5725, B2 => 
                           n6860, ZN => n4400);
   U3220 : NOR2_X1 port map( A1 => n4403, A2 => n4396, ZN => n2480);
   U3221 : NOR2_X1 port map( A1 => n4403, A2 => n4404, ZN => n2479);
   U3222 : AOI22_X1 port map( A1 => n5723, A2 => n2130, B1 => n5720, B2 => 
                           n6743, ZN => n4399);
   U3223 : NOR2_X1 port map( A1 => n4397, A2 => n4379, ZN => n2482);
   U3224 : NOR2_X1 port map( A1 => n4402, A2 => n4383, ZN => n2481);
   U3225 : AOI22_X1 port map( A1 => n5717, A2 => n609, B1 => n5714, B2 => n449,
                           ZN => n4398);
   U3226 : NOR2_X1 port map( A1 => n4405, A2 => n4379, ZN => n2484);
   U3227 : NOR2_X1 port map( A1 => n4405, A2 => n4395, ZN => n2483);
   U3228 : NOR4_X1 port map( A1 => n4406, A2 => n4407, A3 => n4408, A4 => n4409
                           , ZN => n4372);
   U3229 : NAND2_X1 port map( A1 => n4410, A2 => n4411, ZN => n4409);
   U3230 : AOI22_X1 port map( A1 => n5711, A2 => n385, B1 => n5708, B2 => n7052
                           , ZN => n4411);
   U3231 : NOR2_X1 port map( A1 => n4405, A2 => n4403, ZN => n2492);
   U3232 : NOR2_X1 port map( A1 => n4402, A2 => n4403, ZN => n2491);
   U3233 : AOI22_X1 port map( A1 => n5705, A2 => n6827, B1 => n5934, B2 => 
                           OUT1_0_port, ZN => n4410);
   U3234 : NOR2_X1 port map( A1 => n4403, A2 => n4397, ZN => n2493);
   U3235 : NAND2_X1 port map( A1 => n4412, A2 => n4413, ZN => n4408);
   U3236 : AOI22_X1 port map( A1 => n2496, A2 => n417, B1 => n5697, B2 => n6970
                           , ZN => n4413);
   U3237 : NOR2_X1 port map( A1 => n4383, A2 => n4404, ZN => n2497);
   U3238 : NOR2_X1 port map( A1 => n4397, A2 => n4395, ZN => n2496);
   U3239 : NAND2_X1 port map( A1 => n4414, A2 => ADD_RD1(3), ZN => n4397);
   U3240 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => n6054, ZN => n4414);
   U3241 : AOI22_X1 port map( A1 => n5696, A2 => n6795, B1 => n5693, B2 => n545
                           , ZN => n4412);
   U3242 : NOR2_X1 port map( A1 => n4402, A2 => n4395, ZN => n2499);
   U3243 : NAND2_X1 port map( A1 => n4415, A2 => ADD_RD1(3), ZN => n4402);
   U3244 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(0), ZN => n4415);
   U3245 : NOR2_X1 port map( A1 => n4379, A2 => n4404, ZN => n2498);
   U3246 : NAND2_X1 port map( A1 => n4416, A2 => n4417, ZN => n4407);
   U3247 : AOI22_X1 port map( A1 => n5690, A2 => n673, B1 => n5687, B2 => n641,
                           ZN => n4417);
   U3248 : NOR2_X1 port map( A1 => n4396, A2 => n4383, ZN => n2503);
   U3249 : NOR2_X1 port map( A1 => n4395, A2 => n4380, ZN => n2502);
   U3250 : NAND2_X1 port map( A1 => n4418, A2 => n4419, ZN => n4395);
   U3251 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), ZN => n4418);
   U3252 : AOI22_X1 port map( A1 => n5684, A2 => n705, B1 => n5681, B2 => n577,
                           ZN => n4416);
   U3253 : NOR2_X1 port map( A1 => n4405, A2 => n4383, ZN => n2505);
   U3254 : OR2_X1 port map( A1 => n4420, A2 => n6054, ZN => n4405);
   U3255 : OR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n4420);
   U3256 : NOR2_X1 port map( A1 => n4403, A2 => n4380, ZN => n2504);
   U3257 : OR2_X1 port map( A1 => n4421, A2 => n6051, ZN => n4380);
   U3258 : OR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(0), ZN => n4421);
   U3259 : NAND2_X1 port map( A1 => n4422, A2 => n4423, ZN => n4406);
   U3260 : AOI22_X1 port map( A1 => n2508, A2 => n481, B1 => n5673, B2 => n353,
                           ZN => n4423);
   U3261 : NOR2_X1 port map( A1 => n4394, A2 => n4379, ZN => n2509);
   U3262 : NOR2_X1 port map( A1 => n4394, A2 => n4383, ZN => n2508);
   U3263 : NAND2_X1 port map( A1 => n4424, A2 => n4419, ZN => n4383);
   U3264 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n6053, ZN => n4424);
   U3265 : NAND2_X1 port map( A1 => n4425, A2 => ADD_RD1(3), ZN => n4394);
   U3266 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => n6051, ZN => n4425);
   U3267 : AOI22_X1 port map( A1 => n5672, A2 => n513, B1 => n5669, B2 => n321,
                           ZN => n4422);
   U3268 : NOR2_X1 port map( A1 => n4396, A2 => n4379, ZN => n2511);
   U3269 : NAND2_X1 port map( A1 => n4426, A2 => n4419, ZN => n4379);
   U3270 : NOR2_X1 port map( A1 => n6052, A2 => n6053, ZN => n4426);
   U3271 : NAND2_X1 port map( A1 => n4427, A2 => ADD_RD1(3), ZN => n4396);
   U3272 : NOR2_X1 port map( A1 => n6051, A2 => n6054, ZN => n4427);
   U3273 : NOR2_X1 port map( A1 => n4403, A2 => n4381, ZN => n2510);
   U3274 : OR2_X1 port map( A1 => n4428, A2 => n6054, ZN => n4381);
   U3275 : OR2_X1 port map( A1 => ADD_RD1(3), A2 => n6051, ZN => n4428);
   U3276 : NAND2_X1 port map( A1 => n4429, A2 => n4419, ZN => n4403);
   U3277 : NOR2_X1 port map( A1 => n4389, A2 => n4430, ZN => n4419);
   U3280 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD1(3), Z => n4386);
   U3281 : XOR2_X1 port map( A => ADD_RD1(1), B => ADD_WR(1), Z => n4387);
   U3283 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD1(4), Z => n4390);
   U3284 : XOR2_X1 port map( A => ADD_RD1(0), B => ADD_WR(0), Z => n4388);
   U3285 : XOR2_X1 port map( A => ADD_RD1(2), B => ADD_WR(2), Z => n4391);
   U3286 : NAND2_X1 port map( A1 => n4433, A2 => RD1, ZN => n4389);
   U3287 : NOR2_X1 port map( A1 => n4434, A2 => n5932, ZN => n4433);
   U3288 : NOR3_X1 port map( A1 => n4404, A2 => ADD_RD1(2), A3 => ADD_RD1(1), 
                           ZN => n4434);
   U3289 : NAND2_X1 port map( A1 => n4435, A2 => n6054, ZN => n4404);
   U3290 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n4435);
   U3291 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n6052, ZN => n4429);
   U3292 : NAND2_X1 port map( A1 => n4436, A2 => n4437, ZN => n3197);
   U3293 : NOR4_X1 port map( A1 => n4438, A2 => n4439, A3 => n4440, A4 => n4441
                           , ZN => n4437);
   U3294 : OAI21_X1 port map( B1 => n1423, B2 => n5666, A => n4443, ZN => n4441
                           );
   U3295 : NAND2_X1 port map( A1 => n5663, A2 => n6859, ZN => n4443);
   U3296 : OAI21_X1 port map( B1 => n6059, B2 => n5660, A => n4446, ZN => n4440
                           );
   U3297 : AOI22_X1 port map( A1 => n5657, A2 => n6707, B1 => n5654, B2 => 
                           n6987, ZN => n4446);
   U3298 : NAND2_X1 port map( A1 => n4449, A2 => n4450, ZN => n4439);
   U3299 : AOI22_X1 port map( A1 => n5649, A2 => n2830, B1 => n5648, B2 => 
                           n6938, ZN => n4450);
   U3300 : AOI22_X1 port map( A1 => n5645, A2 => n6604, B1 => n5642, B2 => 
                           n6742, ZN => n4449);
   U3302 : AOI22_X1 port map( A1 => n5639, A2 => n2382, B1 => n5636, B2 => 
                           n7019, ZN => n4458);
   U3303 : AOI22_X1 port map( A1 => n5633, A2 => n6667, B1 => n4462, B2 => 
                           n6937, ZN => n4457);
   U3304 : AOI22_X1 port map( A1 => n5627, A2 => n6710, B1 => n5624, B2 => 
                           n7051, ZN => n4456);
   U3305 : AOI22_X1 port map( A1 => n5621, A2 => n640, B1 => n5618, B2 => n480,
                           ZN => n4455);
   U3306 : NOR4_X1 port map( A1 => n4467, A2 => n4468, A3 => n4469, A4 => n4470
                           , ZN => n4436);
   U3307 : NAND2_X1 port map( A1 => n4471, A2 => n4472, ZN => n4470);
   U3308 : AOI22_X1 port map( A1 => n5615, A2 => n416, B1 => n5612, B2 => n7083
                           , ZN => n4472);
   U3309 : AOI22_X1 port map( A1 => n5609, A2 => n6796, B1 => n5935, B2 => 
                           OUT2_31_port, ZN => n4471);
   U3310 : NAND2_X1 port map( A1 => n4476, A2 => n4477, ZN => n4469);
   U3311 : AOI22_X1 port map( A1 => n4478, A2 => n448, B1 => n5601, B2 => n6939
                           , ZN => n4477);
   U3312 : AOI22_X1 port map( A1 => n5600, A2 => n6764, B1 => n5597, B2 => n576
                           , ZN => n4476);
   U3313 : NAND2_X1 port map( A1 => n4482, A2 => n4483, ZN => n4468);
   U3314 : AOI22_X1 port map( A1 => n5594, A2 => n704, B1 => n5591, B2 => n672,
                           ZN => n4483);
   U3315 : AOI22_X1 port map( A1 => n5588, A2 => n736, B1 => n5585, B2 => n608,
                           ZN => n4482);
   U3316 : NAND2_X1 port map( A1 => n4488, A2 => n4489, ZN => n4467);
   U3317 : AOI22_X1 port map( A1 => n4490, A2 => n512, B1 => n5577, B2 => n384,
                           ZN => n4489);
   U3318 : AOI22_X1 port map( A1 => n5576, A2 => n544, B1 => n5573, B2 => n352,
                           ZN => n4488);
   U3319 : NAND2_X1 port map( A1 => n4494, A2 => n4495, ZN => n3196);
   U3320 : NOR4_X1 port map( A1 => n4496, A2 => n4497, A3 => n4498, A4 => n4499
                           , ZN => n4495);
   U3321 : OAI21_X1 port map( B1 => n1424, B2 => n5666, A => n4500, ZN => n4499
                           );
   U3322 : NAND2_X1 port map( A1 => n5663, A2 => n6858, ZN => n4500);
   U3323 : OAI21_X1 port map( B1 => n6060, B2 => n5660, A => n4501, ZN => n4498
                           );
   U3324 : AOI22_X1 port map( A1 => n5657, A2 => n6706, B1 => n5654, B2 => 
                           n6986, ZN => n4501);
   U3325 : NAND2_X1 port map( A1 => n4502, A2 => n4503, ZN => n4497);
   U3326 : AOI22_X1 port map( A1 => n5649, A2 => n2829, B1 => n5648, B2 => 
                           n6936, ZN => n4503);
   U3327 : AOI22_X1 port map( A1 => n5645, A2 => n6605, B1 => n5642, B2 => 
                           n6741, ZN => n4502);
   U3329 : AOI22_X1 port map( A1 => n5639, A2 => n2379, B1 => n5636, B2 => 
                           n7018, ZN => n4507);
   U3330 : AOI22_X1 port map( A1 => n5633, A2 => n6666, B1 => n4462, B2 => 
                           n6935, ZN => n4506);
   U3331 : AOI22_X1 port map( A1 => n5627, A2 => n6709, B1 => n5624, B2 => 
                           n7050, ZN => n4505);
   U3332 : AOI22_X1 port map( A1 => n5621, A2 => n639, B1 => n5618, B2 => n479,
                           ZN => n4504);
   U3333 : NOR4_X1 port map( A1 => n4508, A2 => n4509, A3 => n4510, A4 => n4511
                           , ZN => n4494);
   U3334 : NAND2_X1 port map( A1 => n4512, A2 => n4513, ZN => n4511);
   U3335 : AOI22_X1 port map( A1 => n5615, A2 => n415, B1 => n5612, B2 => n7082
                           , ZN => n4513);
   U3336 : AOI22_X1 port map( A1 => n5609, A2 => n6797, B1 => n5934, B2 => 
                           OUT2_30_port, ZN => n4512);
   U3337 : NAND2_X1 port map( A1 => n4514, A2 => n4515, ZN => n4510);
   U3338 : AOI22_X1 port map( A1 => n4478, A2 => n447, B1 => n5601, B2 => n6940
                           , ZN => n4515);
   U3339 : AOI22_X1 port map( A1 => n5600, A2 => n6765, B1 => n5597, B2 => n575
                           , ZN => n4514);
   U3340 : NAND2_X1 port map( A1 => n4516, A2 => n4517, ZN => n4509);
   U3341 : AOI22_X1 port map( A1 => n5594, A2 => n703, B1 => n5591, B2 => n671,
                           ZN => n4517);
   U3342 : AOI22_X1 port map( A1 => n5588, A2 => n735, B1 => n5585, B2 => n607,
                           ZN => n4516);
   U3343 : NAND2_X1 port map( A1 => n4518, A2 => n4519, ZN => n4508);
   U3344 : AOI22_X1 port map( A1 => n4490, A2 => n511, B1 => n5577, B2 => n383,
                           ZN => n4519);
   U3345 : AOI22_X1 port map( A1 => n5576, A2 => n543, B1 => n5573, B2 => n351,
                           ZN => n4518);
   U3346 : NAND2_X1 port map( A1 => n4520, A2 => n4521, ZN => n3195);
   U3347 : NOR4_X1 port map( A1 => n4522, A2 => n4523, A3 => n4524, A4 => n4525
                           , ZN => n4521);
   U3348 : OAI21_X1 port map( B1 => n1425, B2 => n5666, A => n4526, ZN => n4525
                           );
   U3349 : NAND2_X1 port map( A1 => n5663, A2 => n6857, ZN => n4526);
   U3350 : OAI21_X1 port map( B1 => n6061, B2 => n5660, A => n4527, ZN => n4524
                           );
   U3351 : AOI22_X1 port map( A1 => n5657, A2 => n6705, B1 => n5654, B2 => 
                           n6985, ZN => n4527);
   U3352 : NAND2_X1 port map( A1 => n4528, A2 => n4529, ZN => n4523);
   U3353 : AOI22_X1 port map( A1 => n5649, A2 => n2828, B1 => n5648, B2 => 
                           n6934, ZN => n4529);
   U3354 : AOI22_X1 port map( A1 => n5645, A2 => n6606, B1 => n5642, B2 => 
                           n6740, ZN => n4528);
   U3356 : AOI22_X1 port map( A1 => n5639, A2 => n2376, B1 => n5636, B2 => 
                           n7017, ZN => n4533);
   U3357 : AOI22_X1 port map( A1 => n5633, A2 => n6665, B1 => n4462, B2 => 
                           n6933, ZN => n4532);
   U3358 : AOI22_X1 port map( A1 => n5627, A2 => n6708, B1 => n5624, B2 => 
                           n7049, ZN => n4531);
   U3359 : AOI22_X1 port map( A1 => n5621, A2 => n638, B1 => n5618, B2 => n478,
                           ZN => n4530);
   U3360 : NOR4_X1 port map( A1 => n4534, A2 => n4535, A3 => n4536, A4 => n4537
                           , ZN => n4520);
   U3361 : NAND2_X1 port map( A1 => n4538, A2 => n4539, ZN => n4537);
   U3362 : AOI22_X1 port map( A1 => n5615, A2 => n414, B1 => n5612, B2 => n7081
                           , ZN => n4539);
   U3363 : AOI22_X1 port map( A1 => n5609, A2 => n6798, B1 => n5935, B2 => 
                           OUT2_29_port, ZN => n4538);
   U3364 : NAND2_X1 port map( A1 => n4540, A2 => n4541, ZN => n4536);
   U3365 : AOI22_X1 port map( A1 => n4478, A2 => n446, B1 => n5601, B2 => n6941
                           , ZN => n4541);
   U3366 : AOI22_X1 port map( A1 => n5600, A2 => n6766, B1 => n5597, B2 => n574
                           , ZN => n4540);
   U3367 : NAND2_X1 port map( A1 => n4542, A2 => n4543, ZN => n4535);
   U3368 : AOI22_X1 port map( A1 => n5594, A2 => n702, B1 => n5591, B2 => n670,
                           ZN => n4543);
   U3369 : AOI22_X1 port map( A1 => n5588, A2 => n734, B1 => n5585, B2 => n606,
                           ZN => n4542);
   U3370 : NAND2_X1 port map( A1 => n4544, A2 => n4545, ZN => n4534);
   U3371 : AOI22_X1 port map( A1 => n4490, A2 => n510, B1 => n5577, B2 => n382,
                           ZN => n4545);
   U3372 : AOI22_X1 port map( A1 => n5576, A2 => n542, B1 => n5573, B2 => n350,
                           ZN => n4544);
   U3373 : NAND2_X1 port map( A1 => n4546, A2 => n4547, ZN => n3194);
   U3374 : NOR4_X1 port map( A1 => n4548, A2 => n4549, A3 => n4550, A4 => n4551
                           , ZN => n4547);
   U3375 : OAI21_X1 port map( B1 => n1426, B2 => n5666, A => n4552, ZN => n4551
                           );
   U3376 : NAND2_X1 port map( A1 => n5663, A2 => n6856, ZN => n4552);
   U3377 : OAI21_X1 port map( B1 => n6062, B2 => n5660, A => n4553, ZN => n4550
                           );
   U3378 : AOI22_X1 port map( A1 => n5657, A2 => n6704, B1 => n5654, B2 => 
                           n6984, ZN => n4553);
   U3379 : NAND2_X1 port map( A1 => n4554, A2 => n4555, ZN => n4549);
   U3380 : AOI22_X1 port map( A1 => n5649, A2 => n2827, B1 => n5648, B2 => 
                           n6932, ZN => n4555);
   U3381 : AOI22_X1 port map( A1 => n5645, A2 => n6607, B1 => n5642, B2 => 
                           n6739, ZN => n4554);
   U3383 : AOI22_X1 port map( A1 => n5639, A2 => n2373, B1 => n5636, B2 => 
                           n7016, ZN => n4559);
   U3384 : AOI22_X1 port map( A1 => n5633, A2 => n6664, B1 => n4462, B2 => 
                           n6931, ZN => n4558);
   U3385 : AOI22_X1 port map( A1 => n5627, A2 => n2270, B1 => n5624, B2 => 
                           n7048, ZN => n4557);
   U3386 : AOI22_X1 port map( A1 => n5621, A2 => n637, B1 => n5618, B2 => n477,
                           ZN => n4556);
   U3387 : NOR4_X1 port map( A1 => n4560, A2 => n4561, A3 => n4562, A4 => n4563
                           , ZN => n4546);
   U3388 : NAND2_X1 port map( A1 => n4564, A2 => n4565, ZN => n4563);
   U3389 : AOI22_X1 port map( A1 => n5615, A2 => n413, B1 => n5612, B2 => n7080
                           , ZN => n4565);
   U3390 : AOI22_X1 port map( A1 => n5609, A2 => n6799, B1 => n5934, B2 => 
                           OUT2_28_port, ZN => n4564);
   U3391 : NAND2_X1 port map( A1 => n4566, A2 => n4567, ZN => n4562);
   U3392 : AOI22_X1 port map( A1 => n4478, A2 => n445, B1 => n5601, B2 => n6942
                           , ZN => n4567);
   U3393 : AOI22_X1 port map( A1 => n5600, A2 => n6767, B1 => n5597, B2 => n573
                           , ZN => n4566);
   U3394 : NAND2_X1 port map( A1 => n4568, A2 => n4569, ZN => n4561);
   U3395 : AOI22_X1 port map( A1 => n5594, A2 => n701, B1 => n5591, B2 => n669,
                           ZN => n4569);
   U3396 : AOI22_X1 port map( A1 => n5588, A2 => n733, B1 => n5585, B2 => n605,
                           ZN => n4568);
   U3397 : NAND2_X1 port map( A1 => n4570, A2 => n4571, ZN => n4560);
   U3398 : AOI22_X1 port map( A1 => n4490, A2 => n509, B1 => n5577, B2 => n381,
                           ZN => n4571);
   U3399 : AOI22_X1 port map( A1 => n5576, A2 => n541, B1 => n5573, B2 => n349,
                           ZN => n4570);
   U3400 : NAND2_X1 port map( A1 => n4572, A2 => n4573, ZN => n3193);
   U3401 : NOR4_X1 port map( A1 => n4574, A2 => n4575, A3 => n4576, A4 => n4577
                           , ZN => n4573);
   U3402 : OAI21_X1 port map( B1 => n1427, B2 => n5666, A => n4578, ZN => n4577
                           );
   U3403 : NAND2_X1 port map( A1 => n5663, A2 => n6855, ZN => n4578);
   U3404 : OAI21_X1 port map( B1 => n6063, B2 => n5660, A => n4579, ZN => n4576
                           );
   U3405 : AOI22_X1 port map( A1 => n5657, A2 => n6703, B1 => n5654, B2 => 
                           n6983, ZN => n4579);
   U3406 : NAND2_X1 port map( A1 => n4580, A2 => n4581, ZN => n4575);
   U3407 : AOI22_X1 port map( A1 => n5649, A2 => n2826, B1 => n5648, B2 => 
                           n6930, ZN => n4581);
   U3408 : AOI22_X1 port map( A1 => n5645, A2 => n6608, B1 => n5642, B2 => 
                           n6738, ZN => n4580);
   U3410 : AOI22_X1 port map( A1 => n5639, A2 => n2370, B1 => n5636, B2 => 
                           n7015, ZN => n4585);
   U3411 : AOI22_X1 port map( A1 => n5633, A2 => n6663, B1 => n4462, B2 => 
                           n6929, ZN => n4584);
   U3412 : AOI22_X1 port map( A1 => n5627, A2 => n2265, B1 => n5624, B2 => 
                           n7047, ZN => n4583);
   U3413 : AOI22_X1 port map( A1 => n5621, A2 => n636, B1 => n5618, B2 => n476,
                           ZN => n4582);
   U3414 : NOR4_X1 port map( A1 => n4586, A2 => n4587, A3 => n4588, A4 => n4589
                           , ZN => n4572);
   U3415 : NAND2_X1 port map( A1 => n4590, A2 => n4591, ZN => n4589);
   U3416 : AOI22_X1 port map( A1 => n5615, A2 => n412, B1 => n5612, B2 => n7079
                           , ZN => n4591);
   U3417 : AOI22_X1 port map( A1 => n5609, A2 => n6800, B1 => n5935, B2 => 
                           OUT2_27_port, ZN => n4590);
   U3418 : NAND2_X1 port map( A1 => n4592, A2 => n4593, ZN => n4588);
   U3419 : AOI22_X1 port map( A1 => n5605, A2 => n444, B1 => n5601, B2 => n6943
                           , ZN => n4593);
   U3420 : AOI22_X1 port map( A1 => n5600, A2 => n6768, B1 => n5597, B2 => n572
                           , ZN => n4592);
   U3421 : NAND2_X1 port map( A1 => n4594, A2 => n4595, ZN => n4587);
   U3422 : AOI22_X1 port map( A1 => n5594, A2 => n700, B1 => n5591, B2 => n668,
                           ZN => n4595);
   U3423 : AOI22_X1 port map( A1 => n5588, A2 => n732, B1 => n5585, B2 => n604,
                           ZN => n4594);
   U3424 : NAND2_X1 port map( A1 => n4596, A2 => n4597, ZN => n4586);
   U3425 : AOI22_X1 port map( A1 => n5581, A2 => n508, B1 => n5577, B2 => n380,
                           ZN => n4597);
   U3426 : AOI22_X1 port map( A1 => n5576, A2 => n540, B1 => n5573, B2 => n348,
                           ZN => n4596);
   U3427 : NAND2_X1 port map( A1 => n4598, A2 => n4599, ZN => n3192);
   U3428 : NOR4_X1 port map( A1 => n4600, A2 => n4601, A3 => n4602, A4 => n4603
                           , ZN => n4599);
   U3429 : OAI21_X1 port map( B1 => n1428, B2 => n5666, A => n4604, ZN => n4603
                           );
   U3430 : NAND2_X1 port map( A1 => n5663, A2 => n6854, ZN => n4604);
   U3431 : OAI21_X1 port map( B1 => n6064, B2 => n5660, A => n4605, ZN => n4602
                           );
   U3432 : AOI22_X1 port map( A1 => n5657, A2 => n6702, B1 => n5654, B2 => 
                           n6982, ZN => n4605);
   U3433 : NAND2_X1 port map( A1 => n4606, A2 => n4607, ZN => n4601);
   U3434 : AOI22_X1 port map( A1 => n5649, A2 => n2825, B1 => n5648, B2 => 
                           n6928, ZN => n4607);
   U3435 : AOI22_X1 port map( A1 => n5645, A2 => n6609, B1 => n5642, B2 => 
                           n6737, ZN => n4606);
   U3437 : AOI22_X1 port map( A1 => n5639, A2 => n2367, B1 => n5636, B2 => 
                           n7014, ZN => n4611);
   U3438 : AOI22_X1 port map( A1 => n5633, A2 => n6662, B1 => n4462, B2 => 
                           n6927, ZN => n4610);
   U3439 : AOI22_X1 port map( A1 => n5627, A2 => n2260, B1 => n5624, B2 => 
                           n7046, ZN => n4609);
   U3440 : AOI22_X1 port map( A1 => n5621, A2 => n635, B1 => n5618, B2 => n475,
                           ZN => n4608);
   U3441 : NOR4_X1 port map( A1 => n4612, A2 => n4613, A3 => n4614, A4 => n4615
                           , ZN => n4598);
   U3442 : NAND2_X1 port map( A1 => n4616, A2 => n4617, ZN => n4615);
   U3443 : AOI22_X1 port map( A1 => n5615, A2 => n411, B1 => n5612, B2 => n7078
                           , ZN => n4617);
   U3444 : AOI22_X1 port map( A1 => n5609, A2 => n6801, B1 => n5934, B2 => 
                           OUT2_26_port, ZN => n4616);
   U3445 : NAND2_X1 port map( A1 => n4618, A2 => n4619, ZN => n4614);
   U3446 : AOI22_X1 port map( A1 => n5605, A2 => n443, B1 => n5601, B2 => n6944
                           , ZN => n4619);
   U3447 : AOI22_X1 port map( A1 => n5600, A2 => n6769, B1 => n5597, B2 => n571
                           , ZN => n4618);
   U3448 : NAND2_X1 port map( A1 => n4620, A2 => n4621, ZN => n4613);
   U3449 : AOI22_X1 port map( A1 => n5594, A2 => n699, B1 => n5591, B2 => n667,
                           ZN => n4621);
   U3450 : AOI22_X1 port map( A1 => n5588, A2 => n731, B1 => n5585, B2 => n603,
                           ZN => n4620);
   U3451 : NAND2_X1 port map( A1 => n4622, A2 => n4623, ZN => n4612);
   U3452 : AOI22_X1 port map( A1 => n5581, A2 => n507, B1 => n5577, B2 => n379,
                           ZN => n4623);
   U3453 : AOI22_X1 port map( A1 => n5576, A2 => n539, B1 => n5573, B2 => n347,
                           ZN => n4622);
   U3454 : NAND2_X1 port map( A1 => n4624, A2 => n4625, ZN => n3191);
   U3455 : NOR4_X1 port map( A1 => n4626, A2 => n4627, A3 => n4628, A4 => n4629
                           , ZN => n4625);
   U3456 : OAI21_X1 port map( B1 => n1429, B2 => n5666, A => n4630, ZN => n4629
                           );
   U3457 : NAND2_X1 port map( A1 => n5663, A2 => n6853, ZN => n4630);
   U3458 : OAI21_X1 port map( B1 => n6065, B2 => n5660, A => n4631, ZN => n4628
                           );
   U3459 : AOI22_X1 port map( A1 => n5657, A2 => n6701, B1 => n5654, B2 => 
                           n6981, ZN => n4631);
   U3460 : NAND2_X1 port map( A1 => n4632, A2 => n4633, ZN => n4627);
   U3461 : AOI22_X1 port map( A1 => n5649, A2 => n2824, B1 => n5648, B2 => 
                           n6926, ZN => n4633);
   U3462 : AOI22_X1 port map( A1 => n5645, A2 => n6610, B1 => n5642, B2 => 
                           n6736, ZN => n4632);
   U3464 : AOI22_X1 port map( A1 => n5639, A2 => n2364, B1 => n5636, B2 => 
                           n7013, ZN => n4637);
   U3465 : AOI22_X1 port map( A1 => n5633, A2 => n6661, B1 => n4462, B2 => 
                           n6925, ZN => n4636);
   U3466 : AOI22_X1 port map( A1 => n5627, A2 => n2255, B1 => n5624, B2 => 
                           n7045, ZN => n4635);
   U3467 : AOI22_X1 port map( A1 => n5621, A2 => n634, B1 => n5618, B2 => n474,
                           ZN => n4634);
   U3468 : NOR4_X1 port map( A1 => n4638, A2 => n4639, A3 => n4640, A4 => n4641
                           , ZN => n4624);
   U3469 : NAND2_X1 port map( A1 => n4642, A2 => n4643, ZN => n4641);
   U3470 : AOI22_X1 port map( A1 => n5615, A2 => n410, B1 => n5612, B2 => n7077
                           , ZN => n4643);
   U3471 : AOI22_X1 port map( A1 => n5609, A2 => n6802, B1 => n5935, B2 => 
                           OUT2_25_port, ZN => n4642);
   U3472 : NAND2_X1 port map( A1 => n4644, A2 => n4645, ZN => n4640);
   U3473 : AOI22_X1 port map( A1 => n4478, A2 => n442, B1 => n4479, B2 => n6945
                           , ZN => n4645);
   U3474 : AOI22_X1 port map( A1 => n5600, A2 => n6770, B1 => n5597, B2 => n570
                           , ZN => n4644);
   U3475 : NAND2_X1 port map( A1 => n4646, A2 => n4647, ZN => n4639);
   U3476 : AOI22_X1 port map( A1 => n5594, A2 => n698, B1 => n5591, B2 => n666,
                           ZN => n4647);
   U3477 : AOI22_X1 port map( A1 => n5588, A2 => n730, B1 => n5585, B2 => n602,
                           ZN => n4646);
   U3478 : NAND2_X1 port map( A1 => n4648, A2 => n4649, ZN => n4638);
   U3479 : AOI22_X1 port map( A1 => n4490, A2 => n506, B1 => n4491, B2 => n378,
                           ZN => n4649);
   U3480 : AOI22_X1 port map( A1 => n5576, A2 => n538, B1 => n5573, B2 => n346,
                           ZN => n4648);
   U3481 : NAND2_X1 port map( A1 => n4650, A2 => n4651, ZN => n3190);
   U3482 : NOR4_X1 port map( A1 => n4652, A2 => n4653, A3 => n4654, A4 => n4655
                           , ZN => n4651);
   U3483 : OAI21_X1 port map( B1 => n1430, B2 => n5666, A => n4656, ZN => n4655
                           );
   U3484 : NAND2_X1 port map( A1 => n5663, A2 => n6852, ZN => n4656);
   U3485 : OAI21_X1 port map( B1 => n6066, B2 => n5660, A => n4657, ZN => n4654
                           );
   U3486 : AOI22_X1 port map( A1 => n5657, A2 => n6700, B1 => n5654, B2 => 
                           n6980, ZN => n4657);
   U3487 : NAND2_X1 port map( A1 => n4658, A2 => n4659, ZN => n4653);
   U3488 : AOI22_X1 port map( A1 => n4451, A2 => n2823, B1 => n5648, B2 => 
                           n6924, ZN => n4659);
   U3489 : AOI22_X1 port map( A1 => n5645, A2 => n6611, B1 => n5642, B2 => 
                           n6735, ZN => n4658);
   U3491 : AOI22_X1 port map( A1 => n5639, A2 => n2361, B1 => n5636, B2 => 
                           n7012, ZN => n4663);
   U3492 : AOI22_X1 port map( A1 => n5633, A2 => n6660, B1 => n5629, B2 => 
                           n6923, ZN => n4662);
   U3493 : AOI22_X1 port map( A1 => n5627, A2 => n2250, B1 => n5624, B2 => 
                           n7044, ZN => n4661);
   U3494 : AOI22_X1 port map( A1 => n5621, A2 => n633, B1 => n5618, B2 => n473,
                           ZN => n4660);
   U3495 : NOR4_X1 port map( A1 => n4664, A2 => n4665, A3 => n4666, A4 => n4667
                           , ZN => n4650);
   U3496 : NAND2_X1 port map( A1 => n4668, A2 => n4669, ZN => n4667);
   U3497 : AOI22_X1 port map( A1 => n5615, A2 => n409, B1 => n5612, B2 => n7076
                           , ZN => n4669);
   U3498 : AOI22_X1 port map( A1 => n5609, A2 => n6803, B1 => n5934, B2 => 
                           OUT2_24_port, ZN => n4668);
   U3499 : NAND2_X1 port map( A1 => n4670, A2 => n4671, ZN => n4666);
   U3500 : AOI22_X1 port map( A1 => n4478, A2 => n441, B1 => n4479, B2 => n6946
                           , ZN => n4671);
   U3501 : AOI22_X1 port map( A1 => n5600, A2 => n6771, B1 => n5597, B2 => n569
                           , ZN => n4670);
   U3502 : NAND2_X1 port map( A1 => n4672, A2 => n4673, ZN => n4665);
   U3503 : AOI22_X1 port map( A1 => n5594, A2 => n697, B1 => n5591, B2 => n665,
                           ZN => n4673);
   U3504 : AOI22_X1 port map( A1 => n5588, A2 => n729, B1 => n5585, B2 => n601,
                           ZN => n4672);
   U3505 : NAND2_X1 port map( A1 => n4674, A2 => n4675, ZN => n4664);
   U3506 : AOI22_X1 port map( A1 => n4490, A2 => n505, B1 => n4491, B2 => n377,
                           ZN => n4675);
   U3507 : AOI22_X1 port map( A1 => n5576, A2 => n537, B1 => n5573, B2 => n345,
                           ZN => n4674);
   U3508 : NAND2_X1 port map( A1 => n4676, A2 => n4677, ZN => n3189);
   U3509 : NOR4_X1 port map( A1 => n4678, A2 => n4679, A3 => n4680, A4 => n4681
                           , ZN => n4677);
   U3510 : OAI21_X1 port map( B1 => n1431, B2 => n4442, A => n4682, ZN => n4681
                           );
   U3511 : NAND2_X1 port map( A1 => n5663, A2 => n6851, ZN => n4682);
   U3512 : OAI21_X1 port map( B1 => n5481, B2 => n4445, A => n4683, ZN => n4680
                           );
   U3513 : AOI22_X1 port map( A1 => n5657, A2 => n6699, B1 => n4448, B2 => 
                           n6979, ZN => n4683);
   U3514 : NAND2_X1 port map( A1 => n4684, A2 => n4685, ZN => n4679);
   U3515 : AOI22_X1 port map( A1 => n5649, A2 => n2822, B1 => n4452, B2 => 
                           n6922, ZN => n4685);
   U3516 : AOI22_X1 port map( A1 => n4453, A2 => n6612, B1 => n5642, B2 => 
                           n6734, ZN => n4684);
   U3518 : AOI22_X1 port map( A1 => n5639, A2 => n2358, B1 => n4460, B2 => 
                           n7011, ZN => n4689);
   U3519 : AOI22_X1 port map( A1 => n5633, A2 => n6659, B1 => n5629, B2 => 
                           n6921, ZN => n4688);
   U3520 : AOI22_X1 port map( A1 => n4463, A2 => n2245, B1 => n4464, B2 => 
                           n7043, ZN => n4687);
   U3521 : AOI22_X1 port map( A1 => n4465, A2 => n632, B1 => n5618, B2 => n472,
                           ZN => n4686);
   U3522 : NOR4_X1 port map( A1 => n4690, A2 => n4691, A3 => n4692, A4 => n4693
                           , ZN => n4676);
   U3523 : NAND2_X1 port map( A1 => n4694, A2 => n4695, ZN => n4693);
   U3524 : AOI22_X1 port map( A1 => n5615, A2 => n408, B1 => n4474, B2 => n7075
                           , ZN => n4695);
   U3525 : AOI22_X1 port map( A1 => n5609, A2 => n6804, B1 => n5935, B2 => 
                           OUT2_23_port, ZN => n4694);
   U3526 : NAND2_X1 port map( A1 => n4696, A2 => n4697, ZN => n4692);
   U3527 : AOI22_X1 port map( A1 => n5605, A2 => n440, B1 => n4479, B2 => n6947
                           , ZN => n4697);
   U3528 : AOI22_X1 port map( A1 => n5600, A2 => n6772, B1 => n4481, B2 => n568
                           , ZN => n4696);
   U3529 : NAND2_X1 port map( A1 => n4698, A2 => n4699, ZN => n4691);
   U3530 : AOI22_X1 port map( A1 => n5594, A2 => n696, B1 => n4485, B2 => n664,
                           ZN => n4699);
   U3531 : AOI22_X1 port map( A1 => n5588, A2 => n728, B1 => n4487, B2 => n600,
                           ZN => n4698);
   U3532 : NAND2_X1 port map( A1 => n4700, A2 => n4701, ZN => n4690);
   U3533 : AOI22_X1 port map( A1 => n5581, A2 => n504, B1 => n4491, B2 => n376,
                           ZN => n4701);
   U3534 : AOI22_X1 port map( A1 => n5576, A2 => n536, B1 => n4493, B2 => n344,
                           ZN => n4700);
   U3535 : NAND2_X1 port map( A1 => n4702, A2 => n4703, ZN => n3188);
   U3536 : NOR4_X1 port map( A1 => n4704, A2 => n4705, A3 => n4706, A4 => n4707
                           , ZN => n4703);
   U3537 : OAI21_X1 port map( B1 => n1432, B2 => n4442, A => n4708, ZN => n4707
                           );
   U3538 : NAND2_X1 port map( A1 => n5663, A2 => n6850, ZN => n4708);
   U3539 : OAI21_X1 port map( B1 => n6068, B2 => n4445, A => n4709, ZN => n4706
                           );
   U3540 : AOI22_X1 port map( A1 => n4447, A2 => n6698, B1 => n5654, B2 => 
                           n6978, ZN => n4709);
   U3541 : NAND2_X1 port map( A1 => n4710, A2 => n4711, ZN => n4705);
   U3542 : AOI22_X1 port map( A1 => n4451, A2 => n2821, B1 => n5648, B2 => 
                           n6920, ZN => n4711);
   U3543 : AOI22_X1 port map( A1 => n4453, A2 => n6613, B1 => n5642, B2 => 
                           n6733, ZN => n4710);
   U3545 : AOI22_X1 port map( A1 => n5639, A2 => n2355, B1 => n4460, B2 => 
                           n7010, ZN => n4715);
   U3546 : AOI22_X1 port map( A1 => n5633, A2 => n6658, B1 => n5629, B2 => 
                           n6919, ZN => n4714);
   U3547 : AOI22_X1 port map( A1 => n4463, A2 => n2240, B1 => n4464, B2 => 
                           n7042, ZN => n4713);
   U3548 : AOI22_X1 port map( A1 => n4465, A2 => n631, B1 => n5618, B2 => n471,
                           ZN => n4712);
   U3549 : NOR4_X1 port map( A1 => n4716, A2 => n4717, A3 => n4718, A4 => n4719
                           , ZN => n4702);
   U3550 : NAND2_X1 port map( A1 => n4720, A2 => n4721, ZN => n4719);
   U3551 : AOI22_X1 port map( A1 => n4473, A2 => n407, B1 => n4474, B2 => n7074
                           , ZN => n4721);
   U3552 : AOI22_X1 port map( A1 => n5609, A2 => n6805, B1 => n5932, B2 => 
                           OUT2_22_port, ZN => n4720);
   U3553 : NAND2_X1 port map( A1 => n4722, A2 => n4723, ZN => n4718);
   U3554 : AOI22_X1 port map( A1 => n5605, A2 => n439, B1 => n5601, B2 => n6948
                           , ZN => n4723);
   U3555 : AOI22_X1 port map( A1 => n5600, A2 => n6773, B1 => n4481, B2 => n567
                           , ZN => n4722);
   U3556 : NAND2_X1 port map( A1 => n4724, A2 => n4725, ZN => n4717);
   U3557 : AOI22_X1 port map( A1 => n5594, A2 => n695, B1 => n4485, B2 => n663,
                           ZN => n4725);
   U3558 : AOI22_X1 port map( A1 => n5588, A2 => n727, B1 => n4487, B2 => n599,
                           ZN => n4724);
   U3559 : NAND2_X1 port map( A1 => n4726, A2 => n4727, ZN => n4716);
   U3560 : AOI22_X1 port map( A1 => n5581, A2 => n503, B1 => n5577, B2 => n375,
                           ZN => n4727);
   U3561 : AOI22_X1 port map( A1 => n5576, A2 => n535, B1 => n4493, B2 => n343,
                           ZN => n4726);
   U3562 : NAND2_X1 port map( A1 => n4728, A2 => n4729, ZN => n3187);
   U3563 : NOR4_X1 port map( A1 => n4730, A2 => n4731, A3 => n4732, A4 => n4733
                           , ZN => n4729);
   U3564 : OAI21_X1 port map( B1 => n1433, B2 => n4442, A => n4734, ZN => n4733
                           );
   U3565 : NAND2_X1 port map( A1 => n5663, A2 => n6849, ZN => n4734);
   U3566 : OAI21_X1 port map( B1 => n6069, B2 => n4445, A => n4735, ZN => n4732
                           );
   U3567 : AOI22_X1 port map( A1 => n4447, A2 => n6697, B1 => n5654, B2 => 
                           n6977, ZN => n4735);
   U3568 : NAND2_X1 port map( A1 => n4736, A2 => n4737, ZN => n4731);
   U3569 : AOI22_X1 port map( A1 => n4451, A2 => n2820, B1 => n5648, B2 => 
                           n6918, ZN => n4737);
   U3570 : AOI22_X1 port map( A1 => n4453, A2 => n6614, B1 => n5642, B2 => 
                           n6732, ZN => n4736);
   U3572 : AOI22_X1 port map( A1 => n5639, A2 => n2352, B1 => n4460, B2 => 
                           n7009, ZN => n4741);
   U3573 : AOI22_X1 port map( A1 => n5633, A2 => n6657, B1 => n5629, B2 => 
                           n6917, ZN => n4740);
   U3574 : AOI22_X1 port map( A1 => n4463, A2 => n2235, B1 => n4464, B2 => 
                           n7041, ZN => n4739);
   U3575 : AOI22_X1 port map( A1 => n4465, A2 => n630, B1 => n5618, B2 => n470,
                           ZN => n4738);
   U3576 : NOR4_X1 port map( A1 => n4742, A2 => n4743, A3 => n4744, A4 => n4745
                           , ZN => n4728);
   U3577 : NAND2_X1 port map( A1 => n4746, A2 => n4747, ZN => n4745);
   U3578 : AOI22_X1 port map( A1 => n4473, A2 => n406, B1 => n4474, B2 => n7073
                           , ZN => n4747);
   U3579 : AOI22_X1 port map( A1 => n5609, A2 => n6806, B1 => n5932, B2 => 
                           OUT2_21_port, ZN => n4746);
   U3580 : NAND2_X1 port map( A1 => n4748, A2 => n4749, ZN => n4744);
   U3581 : AOI22_X1 port map( A1 => n5605, A2 => n438, B1 => n4479, B2 => n6949
                           , ZN => n4749);
   U3582 : AOI22_X1 port map( A1 => n5600, A2 => n6774, B1 => n4481, B2 => n566
                           , ZN => n4748);
   U3583 : NAND2_X1 port map( A1 => n4750, A2 => n4751, ZN => n4743);
   U3584 : AOI22_X1 port map( A1 => n5594, A2 => n694, B1 => n4485, B2 => n662,
                           ZN => n4751);
   U3585 : AOI22_X1 port map( A1 => n5588, A2 => n726, B1 => n4487, B2 => n598,
                           ZN => n4750);
   U3586 : NAND2_X1 port map( A1 => n4752, A2 => n4753, ZN => n4742);
   U3587 : AOI22_X1 port map( A1 => n5581, A2 => n502, B1 => n4491, B2 => n374,
                           ZN => n4753);
   U3588 : AOI22_X1 port map( A1 => n5576, A2 => n534, B1 => n4493, B2 => n342,
                           ZN => n4752);
   U3589 : NAND2_X1 port map( A1 => n4754, A2 => n4755, ZN => n3186);
   U3590 : NOR4_X1 port map( A1 => n4756, A2 => n4757, A3 => n4758, A4 => n4759
                           , ZN => n4755);
   U3591 : OAI21_X1 port map( B1 => n1434, B2 => n4442, A => n4760, ZN => n4759
                           );
   U3592 : NAND2_X1 port map( A1 => n5663, A2 => n6848, ZN => n4760);
   U3593 : OAI21_X1 port map( B1 => n6070, B2 => n4445, A => n4761, ZN => n4758
                           );
   U3594 : AOI22_X1 port map( A1 => n4447, A2 => n6696, B1 => n5654, B2 => 
                           n6976, ZN => n4761);
   U3595 : NAND2_X1 port map( A1 => n4762, A2 => n4763, ZN => n4757);
   U3596 : AOI22_X1 port map( A1 => n4451, A2 => n2819, B1 => n5648, B2 => 
                           n6916, ZN => n4763);
   U3597 : AOI22_X1 port map( A1 => n4453, A2 => n6615, B1 => n5642, B2 => 
                           n6731, ZN => n4762);
   U3599 : AOI22_X1 port map( A1 => n5639, A2 => n6763, B1 => n4460, B2 => 
                           n7008, ZN => n4767);
   U3600 : AOI22_X1 port map( A1 => n5633, A2 => n6656, B1 => n5629, B2 => 
                           n6915, ZN => n4766);
   U3601 : AOI22_X1 port map( A1 => n4463, A2 => n2230, B1 => n4464, B2 => 
                           n7040, ZN => n4765);
   U3602 : AOI22_X1 port map( A1 => n4465, A2 => n629, B1 => n5618, B2 => n469,
                           ZN => n4764);
   U3603 : NOR4_X1 port map( A1 => n4768, A2 => n4769, A3 => n4770, A4 => n4771
                           , ZN => n4754);
   U3604 : NAND2_X1 port map( A1 => n4772, A2 => n4773, ZN => n4771);
   U3605 : AOI22_X1 port map( A1 => n4473, A2 => n405, B1 => n4474, B2 => n7072
                           , ZN => n4773);
   U3606 : AOI22_X1 port map( A1 => n5609, A2 => n6807, B1 => n5932, B2 => 
                           OUT2_20_port, ZN => n4772);
   U3607 : NAND2_X1 port map( A1 => n4774, A2 => n4775, ZN => n4770);
   U3608 : AOI22_X1 port map( A1 => n5605, A2 => n437, B1 => n4479, B2 => n6950
                           , ZN => n4775);
   U3609 : AOI22_X1 port map( A1 => n5600, A2 => n6775, B1 => n4481, B2 => n565
                           , ZN => n4774);
   U3610 : NAND2_X1 port map( A1 => n4776, A2 => n4777, ZN => n4769);
   U3611 : AOI22_X1 port map( A1 => n5594, A2 => n693, B1 => n4485, B2 => n661,
                           ZN => n4777);
   U3612 : AOI22_X1 port map( A1 => n5588, A2 => n725, B1 => n4487, B2 => n597,
                           ZN => n4776);
   U3613 : NAND2_X1 port map( A1 => n4778, A2 => n4779, ZN => n4768);
   U3614 : AOI22_X1 port map( A1 => n5581, A2 => n501, B1 => n4491, B2 => n373,
                           ZN => n4779);
   U3615 : AOI22_X1 port map( A1 => n5576, A2 => n533, B1 => n4493, B2 => n341,
                           ZN => n4778);
   U3616 : NAND2_X1 port map( A1 => n4780, A2 => n4781, ZN => n3185);
   U3617 : NOR4_X1 port map( A1 => n4782, A2 => n4783, A3 => n4784, A4 => n4785
                           , ZN => n4781);
   U3618 : OAI21_X1 port map( B1 => n1435, B2 => n4442, A => n4786, ZN => n4785
                           );
   U3619 : NAND2_X1 port map( A1 => n5663, A2 => n6847, ZN => n4786);
   U3620 : OAI21_X1 port map( B1 => n6071, B2 => n4445, A => n4787, ZN => n4784
                           );
   U3621 : AOI22_X1 port map( A1 => n5657, A2 => n6695, B1 => n4448, B2 => 
                           n6975, ZN => n4787);
   U3622 : NAND2_X1 port map( A1 => n4788, A2 => n4789, ZN => n4783);
   U3623 : AOI22_X1 port map( A1 => n4451, A2 => n2818, B1 => n5648, B2 => 
                           n6914, ZN => n4789);
   U3624 : AOI22_X1 port map( A1 => n4453, A2 => n6616, B1 => n5642, B2 => 
                           n6730, ZN => n4788);
   U3626 : AOI22_X1 port map( A1 => n5639, A2 => n6762, B1 => n4460, B2 => 
                           n7007, ZN => n4793);
   U3627 : AOI22_X1 port map( A1 => n5633, A2 => n6655, B1 => n5629, B2 => 
                           n6913, ZN => n4792);
   U3628 : AOI22_X1 port map( A1 => n4463, A2 => n2225, B1 => n4464, B2 => 
                           n7039, ZN => n4791);
   U3629 : AOI22_X1 port map( A1 => n4465, A2 => n628, B1 => n5618, B2 => n468,
                           ZN => n4790);
   U3630 : NOR4_X1 port map( A1 => n4794, A2 => n4795, A3 => n4796, A4 => n4797
                           , ZN => n4780);
   U3631 : NAND2_X1 port map( A1 => n4798, A2 => n4799, ZN => n4797);
   U3632 : AOI22_X1 port map( A1 => n4473, A2 => n404, B1 => n4474, B2 => n7071
                           , ZN => n4799);
   U3633 : AOI22_X1 port map( A1 => n5609, A2 => n6808, B1 => n5932, B2 => 
                           OUT2_19_port, ZN => n4798);
   U3634 : NAND2_X1 port map( A1 => n4800, A2 => n4801, ZN => n4796);
   U3635 : AOI22_X1 port map( A1 => n5605, A2 => n436, B1 => n4479, B2 => n6951
                           , ZN => n4801);
   U3636 : AOI22_X1 port map( A1 => n5600, A2 => n6776, B1 => n4481, B2 => n564
                           , ZN => n4800);
   U3637 : NAND2_X1 port map( A1 => n4802, A2 => n4803, ZN => n4795);
   U3638 : AOI22_X1 port map( A1 => n5594, A2 => n692, B1 => n4485, B2 => n660,
                           ZN => n4803);
   U3639 : AOI22_X1 port map( A1 => n5588, A2 => n724, B1 => n4487, B2 => n596,
                           ZN => n4802);
   U3640 : NAND2_X1 port map( A1 => n4804, A2 => n4805, ZN => n4794);
   U3641 : AOI22_X1 port map( A1 => n5581, A2 => n500, B1 => n4491, B2 => n372,
                           ZN => n4805);
   U3642 : AOI22_X1 port map( A1 => n5576, A2 => n532, B1 => n4493, B2 => n340,
                           ZN => n4804);
   U3643 : NAND2_X1 port map( A1 => n4806, A2 => n4807, ZN => n3184);
   U3644 : NOR4_X1 port map( A1 => n4808, A2 => n4809, A3 => n4810, A4 => n4811
                           , ZN => n4807);
   U3645 : OAI21_X1 port map( B1 => n1436, B2 => n4442, A => n4812, ZN => n4811
                           );
   U3646 : NAND2_X1 port map( A1 => n4444, A2 => n6846, ZN => n4812);
   U3647 : OAI21_X1 port map( B1 => n6072, B2 => n4445, A => n4813, ZN => n4810
                           );
   U3648 : AOI22_X1 port map( A1 => n5657, A2 => n6694, B1 => n4448, B2 => 
                           n6974, ZN => n4813);
   U3649 : NAND2_X1 port map( A1 => n4814, A2 => n4815, ZN => n4809);
   U3650 : AOI22_X1 port map( A1 => n4451, A2 => n2817, B1 => n5648, B2 => 
                           n6912, ZN => n4815);
   U3651 : AOI22_X1 port map( A1 => n5645, A2 => n6617, B1 => n4454, B2 => 
                           n6729, ZN => n4814);
   U3653 : AOI22_X1 port map( A1 => n5639, A2 => n6761, B1 => n5636, B2 => 
                           n7006, ZN => n4819);
   U3654 : AOI22_X1 port map( A1 => n5633, A2 => n6654, B1 => n5629, B2 => 
                           n6911, ZN => n4818);
   U3655 : AOI22_X1 port map( A1 => n5627, A2 => n2220, B1 => n5624, B2 => 
                           n7038, ZN => n4817);
   U3656 : AOI22_X1 port map( A1 => n5621, A2 => n627, B1 => n4466, B2 => n467,
                           ZN => n4816);
   U3657 : NOR4_X1 port map( A1 => n4820, A2 => n4821, A3 => n4822, A4 => n4823
                           , ZN => n4806);
   U3658 : NAND2_X1 port map( A1 => n4824, A2 => n4825, ZN => n4823);
   U3659 : AOI22_X1 port map( A1 => n4473, A2 => n403, B1 => n4474, B2 => n7070
                           , ZN => n4825);
   U3660 : AOI22_X1 port map( A1 => n5609, A2 => n6809, B1 => n5932, B2 => 
                           OUT2_18_port, ZN => n4824);
   U3661 : NAND2_X1 port map( A1 => n4826, A2 => n4827, ZN => n4822);
   U3662 : AOI22_X1 port map( A1 => n5605, A2 => n435, B1 => n4479, B2 => n6952
                           , ZN => n4827);
   U3663 : AOI22_X1 port map( A1 => n5600, A2 => n6777, B1 => n4481, B2 => n563
                           , ZN => n4826);
   U3664 : NAND2_X1 port map( A1 => n4828, A2 => n4829, ZN => n4821);
   U3665 : AOI22_X1 port map( A1 => n5594, A2 => n691, B1 => n4485, B2 => n659,
                           ZN => n4829);
   U3666 : AOI22_X1 port map( A1 => n5588, A2 => n723, B1 => n4487, B2 => n595,
                           ZN => n4828);
   U3667 : NAND2_X1 port map( A1 => n4830, A2 => n4831, ZN => n4820);
   U3668 : AOI22_X1 port map( A1 => n5581, A2 => n499, B1 => n4491, B2 => n371,
                           ZN => n4831);
   U3669 : AOI22_X1 port map( A1 => n5576, A2 => n531, B1 => n4493, B2 => n339,
                           ZN => n4830);
   U3670 : NAND2_X1 port map( A1 => n4832, A2 => n4833, ZN => n3183);
   U3671 : NOR4_X1 port map( A1 => n4834, A2 => n4835, A3 => n4836, A4 => n4837
                           , ZN => n4833);
   U3672 : OAI21_X1 port map( B1 => n1437, B2 => n4442, A => n4838, ZN => n4837
                           );
   U3673 : NAND2_X1 port map( A1 => n4444, A2 => n6845, ZN => n4838);
   U3674 : OAI21_X1 port map( B1 => n5499, B2 => n4445, A => n4839, ZN => n4836
                           );
   U3675 : AOI22_X1 port map( A1 => n5657, A2 => n6693, B1 => n4448, B2 => 
                           n6973, ZN => n4839);
   U3676 : NAND2_X1 port map( A1 => n4840, A2 => n4841, ZN => n4835);
   U3677 : AOI22_X1 port map( A1 => n4451, A2 => n2816, B1 => n5648, B2 => 
                           n6910, ZN => n4841);
   U3678 : AOI22_X1 port map( A1 => n5645, A2 => n6618, B1 => n4454, B2 => 
                           n6728, ZN => n4840);
   U3680 : AOI22_X1 port map( A1 => n4459, A2 => n6760, B1 => n5636, B2 => 
                           n7005, ZN => n4845);
   U3681 : AOI22_X1 port map( A1 => n4461, A2 => n6653, B1 => n5629, B2 => 
                           n6909, ZN => n4844);
   U3682 : AOI22_X1 port map( A1 => n5627, A2 => n2215, B1 => n5624, B2 => 
                           n7037, ZN => n4843);
   U3683 : AOI22_X1 port map( A1 => n5621, A2 => n626, B1 => n4466, B2 => n466,
                           ZN => n4842);
   U3684 : NOR4_X1 port map( A1 => n4846, A2 => n4847, A3 => n4848, A4 => n4849
                           , ZN => n4832);
   U3685 : NAND2_X1 port map( A1 => n4850, A2 => n4851, ZN => n4849);
   U3686 : AOI22_X1 port map( A1 => n5615, A2 => n402, B1 => n5612, B2 => n7069
                           , ZN => n4851);
   U3687 : AOI22_X1 port map( A1 => n4475, A2 => n6810, B1 => n5934, B2 => 
                           OUT2_17_port, ZN => n4850);
   U3688 : NAND2_X1 port map( A1 => n4852, A2 => n4853, ZN => n4848);
   U3689 : AOI22_X1 port map( A1 => n5605, A2 => n434, B1 => n4479, B2 => n6953
                           , ZN => n4853);
   U3690 : AOI22_X1 port map( A1 => n4480, A2 => n6778, B1 => n5597, B2 => n562
                           , ZN => n4852);
   U3691 : NAND2_X1 port map( A1 => n4854, A2 => n4855, ZN => n4847);
   U3692 : AOI22_X1 port map( A1 => n5594, A2 => n690, B1 => n5591, B2 => n658,
                           ZN => n4855);
   U3693 : AOI22_X1 port map( A1 => n4486, A2 => n722, B1 => n5585, B2 => n594,
                           ZN => n4854);
   U3694 : NAND2_X1 port map( A1 => n4856, A2 => n4857, ZN => n4846);
   U3695 : AOI22_X1 port map( A1 => n5581, A2 => n498, B1 => n4491, B2 => n370,
                           ZN => n4857);
   U3696 : AOI22_X1 port map( A1 => n4492, A2 => n530, B1 => n5573, B2 => n338,
                           ZN => n4856);
   U3697 : NAND2_X1 port map( A1 => n4858, A2 => n4859, ZN => n3182);
   U3698 : NOR4_X1 port map( A1 => n4860, A2 => n4861, A3 => n4862, A4 => n4863
                           , ZN => n4859);
   U3699 : OAI21_X1 port map( B1 => n1438, B2 => n4442, A => n4864, ZN => n4863
                           );
   U3700 : NAND2_X1 port map( A1 => n4444, A2 => n6844, ZN => n4864);
   U3701 : OAI21_X1 port map( B1 => n6074, B2 => n4445, A => n4865, ZN => n4862
                           );
   U3702 : AOI22_X1 port map( A1 => n5657, A2 => n6692, B1 => n4448, B2 => 
                           n6972, ZN => n4865);
   U3703 : NAND2_X1 port map( A1 => n4866, A2 => n4867, ZN => n4861);
   U3704 : AOI22_X1 port map( A1 => n4451, A2 => n2815, B1 => n4452, B2 => 
                           n6908, ZN => n4867);
   U3705 : AOI22_X1 port map( A1 => n5645, A2 => n6619, B1 => n4454, B2 => 
                           n6727, ZN => n4866);
   U3707 : AOI22_X1 port map( A1 => n4459, A2 => n6759, B1 => n5636, B2 => 
                           n7004, ZN => n4871);
   U3708 : AOI22_X1 port map( A1 => n4461, A2 => n6652, B1 => n5629, B2 => 
                           n6907, ZN => n4870);
   U3709 : AOI22_X1 port map( A1 => n5627, A2 => n2210, B1 => n5624, B2 => 
                           n7036, ZN => n4869);
   U3710 : AOI22_X1 port map( A1 => n5621, A2 => n625, B1 => n4466, B2 => n465,
                           ZN => n4868);
   U3711 : NOR4_X1 port map( A1 => n4872, A2 => n4873, A3 => n4874, A4 => n4875
                           , ZN => n4858);
   U3712 : NAND2_X1 port map( A1 => n4876, A2 => n4877, ZN => n4875);
   U3713 : AOI22_X1 port map( A1 => n5615, A2 => n401, B1 => n5612, B2 => n7068
                           , ZN => n4877);
   U3714 : AOI22_X1 port map( A1 => n4475, A2 => n6811, B1 => n5932, B2 => 
                           OUT2_16_port, ZN => n4876);
   U3715 : NAND2_X1 port map( A1 => n4878, A2 => n4879, ZN => n4874);
   U3716 : AOI22_X1 port map( A1 => n5605, A2 => n433, B1 => n4479, B2 => n6954
                           , ZN => n4879);
   U3717 : AOI22_X1 port map( A1 => n4480, A2 => n6779, B1 => n5597, B2 => n561
                           , ZN => n4878);
   U3718 : NAND2_X1 port map( A1 => n4880, A2 => n4881, ZN => n4873);
   U3719 : AOI22_X1 port map( A1 => n4484, A2 => n689, B1 => n5591, B2 => n657,
                           ZN => n4881);
   U3720 : AOI22_X1 port map( A1 => n4486, A2 => n721, B1 => n5585, B2 => n593,
                           ZN => n4880);
   U3721 : NAND2_X1 port map( A1 => n4882, A2 => n4883, ZN => n4872);
   U3722 : AOI22_X1 port map( A1 => n5581, A2 => n497, B1 => n4491, B2 => n369,
                           ZN => n4883);
   U3723 : AOI22_X1 port map( A1 => n4492, A2 => n529, B1 => n5573, B2 => n337,
                           ZN => n4882);
   U3724 : NAND2_X1 port map( A1 => n4884, A2 => n4885, ZN => n3181);
   U3725 : NOR4_X1 port map( A1 => n4886, A2 => n4887, A3 => n4888, A4 => n4889
                           , ZN => n4885);
   U3726 : OAI21_X1 port map( B1 => n1439, B2 => n4442, A => n4890, ZN => n4889
                           );
   U3727 : NAND2_X1 port map( A1 => n5663, A2 => n6843, ZN => n4890);
   U3728 : OAI21_X1 port map( B1 => n6075, B2 => n4445, A => n4891, ZN => n4888
                           );
   U3729 : AOI22_X1 port map( A1 => n5657, A2 => n6691, B1 => n5654, B2 => 
                           n6971, ZN => n4891);
   U3730 : NAND2_X1 port map( A1 => n4892, A2 => n4893, ZN => n4887);
   U3731 : AOI22_X1 port map( A1 => n5649, A2 => n2814, B1 => n5648, B2 => 
                           n6906, ZN => n4893);
   U3732 : AOI22_X1 port map( A1 => n5645, A2 => n6620, B1 => n5642, B2 => 
                           n6726, ZN => n4892);
   U3734 : AOI22_X1 port map( A1 => n5639, A2 => n6758, B1 => n5636, B2 => 
                           n7003, ZN => n4897);
   U3735 : AOI22_X1 port map( A1 => n5633, A2 => n6651, B1 => n5629, B2 => 
                           n6905, ZN => n4896);
   U3736 : AOI22_X1 port map( A1 => n5627, A2 => n2205, B1 => n5624, B2 => 
                           n7035, ZN => n4895);
   U3737 : AOI22_X1 port map( A1 => n5621, A2 => n624, B1 => n5618, B2 => n464,
                           ZN => n4894);
   U3738 : NOR4_X1 port map( A1 => n4898, A2 => n4899, A3 => n4900, A4 => n4901
                           , ZN => n4884);
   U3739 : NAND2_X1 port map( A1 => n4902, A2 => n4903, ZN => n4901);
   U3740 : AOI22_X1 port map( A1 => n5615, A2 => n400, B1 => n5612, B2 => n7067
                           , ZN => n4903);
   U3741 : AOI22_X1 port map( A1 => n4475, A2 => n6812, B1 => n5935, B2 => 
                           OUT2_15_port, ZN => n4902);
   U3742 : NAND2_X1 port map( A1 => n4904, A2 => n4905, ZN => n4900);
   U3743 : AOI22_X1 port map( A1 => n5605, A2 => n432, B1 => n4479, B2 => n6955
                           , ZN => n4905);
   U3744 : AOI22_X1 port map( A1 => n4480, A2 => n6780, B1 => n5597, B2 => n560
                           , ZN => n4904);
   U3745 : NAND2_X1 port map( A1 => n4906, A2 => n4907, ZN => n4899);
   U3746 : AOI22_X1 port map( A1 => n4484, A2 => n688, B1 => n5591, B2 => n656,
                           ZN => n4907);
   U3747 : AOI22_X1 port map( A1 => n4486, A2 => n720, B1 => n5585, B2 => n592,
                           ZN => n4906);
   U3748 : NAND2_X1 port map( A1 => n4908, A2 => n4909, ZN => n4898);
   U3749 : AOI22_X1 port map( A1 => n5581, A2 => n496, B1 => n4491, B2 => n368,
                           ZN => n4909);
   U3750 : AOI22_X1 port map( A1 => n4492, A2 => n528, B1 => n5573, B2 => n336,
                           ZN => n4908);
   U3751 : NAND2_X1 port map( A1 => n4910, A2 => n4911, ZN => n3180);
   U3752 : NOR4_X1 port map( A1 => n4912, A2 => n4913, A3 => n4914, A4 => n4915
                           , ZN => n4911);
   U3753 : OAI21_X1 port map( B1 => n1440, B2 => n4442, A => n4916, ZN => n4915
                           );
   U3754 : NAND2_X1 port map( A1 => n4444, A2 => n6842, ZN => n4916);
   U3755 : OAI21_X1 port map( B1 => n6076, B2 => n4445, A => n4917, ZN => n4914
                           );
   U3756 : AOI22_X1 port map( A1 => n5657, A2 => n6690, B1 => n4448, B2 => 
                           n6904, ZN => n4917);
   U3757 : NAND2_X1 port map( A1 => n4918, A2 => n4919, ZN => n4913);
   U3758 : AOI22_X1 port map( A1 => n4451, A2 => n2813, B1 => n4452, B2 => 
                           n6903, ZN => n4919);
   U3759 : AOI22_X1 port map( A1 => n5645, A2 => n6621, B1 => n4454, B2 => 
                           n6725, ZN => n4918);
   U3761 : AOI22_X1 port map( A1 => n4459, A2 => n6757, B1 => n5636, B2 => 
                           n7002, ZN => n4923);
   U3762 : AOI22_X1 port map( A1 => n4461, A2 => n6650, B1 => n5629, B2 => 
                           n6902, ZN => n4922);
   U3763 : AOI22_X1 port map( A1 => n5627, A2 => n2200, B1 => n5624, B2 => 
                           n7034, ZN => n4921);
   U3764 : AOI22_X1 port map( A1 => n5621, A2 => n623, B1 => n4466, B2 => n463,
                           ZN => n4920);
   U3765 : NOR4_X1 port map( A1 => n4924, A2 => n4925, A3 => n4926, A4 => n4927
                           , ZN => n4910);
   U3766 : NAND2_X1 port map( A1 => n4928, A2 => n4929, ZN => n4927);
   U3767 : AOI22_X1 port map( A1 => n5615, A2 => n399, B1 => n5612, B2 => n7066
                           , ZN => n4929);
   U3768 : AOI22_X1 port map( A1 => n4475, A2 => n6813, B1 => n5932, B2 => 
                           OUT2_14_port, ZN => n4928);
   U3769 : NAND2_X1 port map( A1 => n4930, A2 => n4931, ZN => n4926);
   U3770 : AOI22_X1 port map( A1 => n5605, A2 => n431, B1 => n4479, B2 => n6956
                           , ZN => n4931);
   U3771 : AOI22_X1 port map( A1 => n4480, A2 => n6781, B1 => n5597, B2 => n559
                           , ZN => n4930);
   U3772 : NAND2_X1 port map( A1 => n4932, A2 => n4933, ZN => n4925);
   U3773 : AOI22_X1 port map( A1 => n4484, A2 => n687, B1 => n5591, B2 => n655,
                           ZN => n4933);
   U3774 : AOI22_X1 port map( A1 => n4486, A2 => n719, B1 => n5585, B2 => n591,
                           ZN => n4932);
   U3775 : NAND2_X1 port map( A1 => n4934, A2 => n4935, ZN => n4924);
   U3776 : AOI22_X1 port map( A1 => n5581, A2 => n495, B1 => n4491, B2 => n367,
                           ZN => n4935);
   U3777 : AOI22_X1 port map( A1 => n4492, A2 => n527, B1 => n5573, B2 => n335,
                           ZN => n4934);
   U3778 : NAND2_X1 port map( A1 => n4936, A2 => n4937, ZN => n3179);
   U3779 : NOR4_X1 port map( A1 => n4938, A2 => n4939, A3 => n4940, A4 => n4941
                           , ZN => n4937);
   U3780 : OAI21_X1 port map( B1 => n1441, B2 => n4442, A => n4942, ZN => n4941
                           );
   U3781 : NAND2_X1 port map( A1 => n4444, A2 => n6841, ZN => n4942);
   U3782 : OAI21_X1 port map( B1 => n6077, B2 => n4445, A => n4943, ZN => n4940
                           );
   U3783 : AOI22_X1 port map( A1 => n4447, A2 => n6689, B1 => n5654, B2 => 
                           n6901, ZN => n4943);
   U3784 : NAND2_X1 port map( A1 => n4944, A2 => n4945, ZN => n4939);
   U3785 : AOI22_X1 port map( A1 => n4451, A2 => n2812, B1 => n4452, B2 => 
                           n6900, ZN => n4945);
   U3786 : AOI22_X1 port map( A1 => n5645, A2 => n6622, B1 => n4454, B2 => 
                           n6724, ZN => n4944);
   U3788 : AOI22_X1 port map( A1 => n4459, A2 => n6756, B1 => n5636, B2 => 
                           n7001, ZN => n4949);
   U3789 : AOI22_X1 port map( A1 => n4461, A2 => n6649, B1 => n5629, B2 => 
                           n6899, ZN => n4948);
   U3790 : AOI22_X1 port map( A1 => n5627, A2 => n2195, B1 => n5624, B2 => 
                           n7033, ZN => n4947);
   U3791 : AOI22_X1 port map( A1 => n5621, A2 => n622, B1 => n4466, B2 => n462,
                           ZN => n4946);
   U3792 : NOR4_X1 port map( A1 => n4950, A2 => n4951, A3 => n4952, A4 => n4953
                           , ZN => n4936);
   U3793 : NAND2_X1 port map( A1 => n4954, A2 => n4955, ZN => n4953);
   U3794 : AOI22_X1 port map( A1 => n5615, A2 => n398, B1 => n5612, B2 => n7065
                           , ZN => n4955);
   U3795 : AOI22_X1 port map( A1 => n4475, A2 => n6814, B1 => n5932, B2 => 
                           OUT2_13_port, ZN => n4954);
   U3796 : NAND2_X1 port map( A1 => n4956, A2 => n4957, ZN => n4952);
   U3797 : AOI22_X1 port map( A1 => n5605, A2 => n430, B1 => n4479, B2 => n6957
                           , ZN => n4957);
   U3798 : AOI22_X1 port map( A1 => n4480, A2 => n6782, B1 => n5597, B2 => n558
                           , ZN => n4956);
   U3799 : NAND2_X1 port map( A1 => n4958, A2 => n4959, ZN => n4951);
   U3800 : AOI22_X1 port map( A1 => n4484, A2 => n686, B1 => n5591, B2 => n654,
                           ZN => n4959);
   U3801 : AOI22_X1 port map( A1 => n4486, A2 => n718, B1 => n5585, B2 => n590,
                           ZN => n4958);
   U3802 : NAND2_X1 port map( A1 => n4960, A2 => n4961, ZN => n4950);
   U3803 : AOI22_X1 port map( A1 => n5581, A2 => n494, B1 => n4491, B2 => n366,
                           ZN => n4961);
   U3804 : AOI22_X1 port map( A1 => n4492, A2 => n526, B1 => n5573, B2 => n334,
                           ZN => n4960);
   U3805 : NAND2_X1 port map( A1 => n4962, A2 => n4963, ZN => n3178);
   U3806 : NOR4_X1 port map( A1 => n4964, A2 => n4965, A3 => n4966, A4 => n4967
                           , ZN => n4963);
   U3807 : OAI21_X1 port map( B1 => n1442, B2 => n4442, A => n4968, ZN => n4967
                           );
   U3808 : NAND2_X1 port map( A1 => n4444, A2 => n6840, ZN => n4968);
   U3809 : OAI21_X1 port map( B1 => n6078, B2 => n4445, A => n4969, ZN => n4966
                           );
   U3810 : AOI22_X1 port map( A1 => n4447, A2 => n6688, B1 => n5654, B2 => 
                           n6898, ZN => n4969);
   U3811 : NAND2_X1 port map( A1 => n4970, A2 => n4971, ZN => n4965);
   U3812 : AOI22_X1 port map( A1 => n4451, A2 => n2811, B1 => n4452, B2 => 
                           n6897, ZN => n4971);
   U3813 : AOI22_X1 port map( A1 => n5645, A2 => n6623, B1 => n4454, B2 => 
                           n6723, ZN => n4970);
   U3815 : AOI22_X1 port map( A1 => n4459, A2 => n6755, B1 => n5636, B2 => 
                           n7000, ZN => n4975);
   U3816 : AOI22_X1 port map( A1 => n4461, A2 => n6648, B1 => n5629, B2 => 
                           n6896, ZN => n4974);
   U3817 : AOI22_X1 port map( A1 => n5627, A2 => n2190, B1 => n5624, B2 => 
                           n7032, ZN => n4973);
   U3818 : AOI22_X1 port map( A1 => n5621, A2 => n621, B1 => n4466, B2 => n461,
                           ZN => n4972);
   U3819 : NOR4_X1 port map( A1 => n4976, A2 => n4977, A3 => n4978, A4 => n4979
                           , ZN => n4962);
   U3820 : NAND2_X1 port map( A1 => n4980, A2 => n4981, ZN => n4979);
   U3821 : AOI22_X1 port map( A1 => n5615, A2 => n397, B1 => n5612, B2 => n7064
                           , ZN => n4981);
   U3822 : AOI22_X1 port map( A1 => n5609, A2 => n6815, B1 => n5932, B2 => 
                           OUT2_12_port, ZN => n4980);
   U3823 : NAND2_X1 port map( A1 => n4982, A2 => n4983, ZN => n4978);
   U3824 : AOI22_X1 port map( A1 => n5605, A2 => n429, B1 => n5601, B2 => n6958
                           , ZN => n4983);
   U3825 : AOI22_X1 port map( A1 => n5600, A2 => n6783, B1 => n5597, B2 => n557
                           , ZN => n4982);
   U3826 : NAND2_X1 port map( A1 => n4984, A2 => n4985, ZN => n4977);
   U3827 : AOI22_X1 port map( A1 => n5594, A2 => n685, B1 => n5591, B2 => n653,
                           ZN => n4985);
   U3828 : AOI22_X1 port map( A1 => n5588, A2 => n717, B1 => n5585, B2 => n589,
                           ZN => n4984);
   U3829 : NAND2_X1 port map( A1 => n4986, A2 => n4987, ZN => n4976);
   U3830 : AOI22_X1 port map( A1 => n5581, A2 => n493, B1 => n5577, B2 => n365,
                           ZN => n4987);
   U3831 : AOI22_X1 port map( A1 => n5576, A2 => n525, B1 => n5573, B2 => n333,
                           ZN => n4986);
   U3832 : NAND2_X1 port map( A1 => n4988, A2 => n4989, ZN => n3177);
   U3833 : NOR4_X1 port map( A1 => n4990, A2 => n4991, A3 => n4992, A4 => n4993
                           , ZN => n4989);
   U3834 : OAI21_X1 port map( B1 => n1443, B2 => n4442, A => n4994, ZN => n4993
                           );
   U3835 : NAND2_X1 port map( A1 => n4444, A2 => n6839, ZN => n4994);
   U3836 : OAI21_X1 port map( B1 => n6079, B2 => n4445, A => n4995, ZN => n4992
                           );
   U3837 : AOI22_X1 port map( A1 => n4447, A2 => n6687, B1 => n4448, B2 => 
                           n6895, ZN => n4995);
   U3838 : NAND2_X1 port map( A1 => n4996, A2 => n4997, ZN => n4991);
   U3839 : AOI22_X1 port map( A1 => n5649, A2 => n2810, B1 => n4452, B2 => 
                           n6894, ZN => n4997);
   U3840 : AOI22_X1 port map( A1 => n4453, A2 => n6624, B1 => n4454, B2 => 
                           n6722, ZN => n4996);
   U3842 : AOI22_X1 port map( A1 => n4459, A2 => n6754, B1 => n4460, B2 => 
                           n6999, ZN => n5001);
   U3843 : AOI22_X1 port map( A1 => n4461, A2 => n6647, B1 => n5629, B2 => 
                           n6893, ZN => n5000);
   U3844 : AOI22_X1 port map( A1 => n4463, A2 => n2185, B1 => n4464, B2 => 
                           n7031, ZN => n4999);
   U3845 : AOI22_X1 port map( A1 => n4465, A2 => n620, B1 => n4466, B2 => n460,
                           ZN => n4998);
   U3846 : NOR4_X1 port map( A1 => n5002, A2 => n5003, A3 => n5004, A4 => n5005
                           , ZN => n4988);
   U3847 : NAND2_X1 port map( A1 => n5006, A2 => n5007, ZN => n5005);
   U3848 : AOI22_X1 port map( A1 => n4473, A2 => n396, B1 => n4474, B2 => n7063
                           , ZN => n5007);
   U3849 : AOI22_X1 port map( A1 => n4475, A2 => n6816, B1 => n5932, B2 => 
                           OUT2_11_port, ZN => n5006);
   U3850 : NAND2_X1 port map( A1 => n5008, A2 => n5009, ZN => n5004);
   U3851 : AOI22_X1 port map( A1 => n5605, A2 => n428, B1 => n5601, B2 => n6959
                           , ZN => n5009);
   U3852 : AOI22_X1 port map( A1 => n4480, A2 => n6784, B1 => n4481, B2 => n556
                           , ZN => n5008);
   U3853 : NAND2_X1 port map( A1 => n5010, A2 => n5011, ZN => n5003);
   U3854 : AOI22_X1 port map( A1 => n4484, A2 => n684, B1 => n4485, B2 => n652,
                           ZN => n5011);
   U3855 : AOI22_X1 port map( A1 => n4486, A2 => n716, B1 => n4487, B2 => n588,
                           ZN => n5010);
   U3856 : NAND2_X1 port map( A1 => n5012, A2 => n5013, ZN => n5002);
   U3857 : AOI22_X1 port map( A1 => n5581, A2 => n492, B1 => n5577, B2 => n364,
                           ZN => n5013);
   U3858 : AOI22_X1 port map( A1 => n4492, A2 => n524, B1 => n4493, B2 => n332,
                           ZN => n5012);
   U3859 : NAND2_X1 port map( A1 => n5014, A2 => n5015, ZN => n3176);
   U3860 : NOR4_X1 port map( A1 => n5016, A2 => n5017, A3 => n5018, A4 => n5019
                           , ZN => n5015);
   U3861 : OAI21_X1 port map( B1 => n1444, B2 => n4442, A => n5020, ZN => n5019
                           );
   U3862 : NAND2_X1 port map( A1 => n4444, A2 => n6838, ZN => n5020);
   U3863 : OAI21_X1 port map( B1 => n6080, B2 => n4445, A => n5021, ZN => n5018
                           );
   U3864 : AOI22_X1 port map( A1 => n4447, A2 => n6686, B1 => n4448, B2 => 
                           n6892, ZN => n5021);
   U3865 : NAND2_X1 port map( A1 => n5022, A2 => n5023, ZN => n5017);
   U3866 : AOI22_X1 port map( A1 => n5649, A2 => n2809, B1 => n4452, B2 => 
                           n6891, ZN => n5023);
   U3867 : AOI22_X1 port map( A1 => n4453, A2 => n6625, B1 => n4454, B2 => 
                           n6721, ZN => n5022);
   U3869 : AOI22_X1 port map( A1 => n4459, A2 => n6753, B1 => n4460, B2 => 
                           n6998, ZN => n5027);
   U3870 : AOI22_X1 port map( A1 => n4461, A2 => n6646, B1 => n5629, B2 => 
                           n6890, ZN => n5026);
   U3871 : AOI22_X1 port map( A1 => n4463, A2 => n2180, B1 => n4464, B2 => 
                           n7030, ZN => n5025);
   U3872 : AOI22_X1 port map( A1 => n4465, A2 => n619, B1 => n4466, B2 => n459,
                           ZN => n5024);
   U3873 : NOR4_X1 port map( A1 => n5028, A2 => n5029, A3 => n5030, A4 => n5031
                           , ZN => n5014);
   U3874 : NAND2_X1 port map( A1 => n5032, A2 => n5033, ZN => n5031);
   U3875 : AOI22_X1 port map( A1 => n4473, A2 => n395, B1 => n4474, B2 => n7062
                           , ZN => n5033);
   U3876 : AOI22_X1 port map( A1 => n4475, A2 => n6817, B1 => n5935, B2 => 
                           OUT2_10_port, ZN => n5032);
   U3877 : NAND2_X1 port map( A1 => n5034, A2 => n5035, ZN => n5030);
   U3878 : AOI22_X1 port map( A1 => n5605, A2 => n427, B1 => n5601, B2 => n6960
                           , ZN => n5035);
   U3879 : AOI22_X1 port map( A1 => n4480, A2 => n6785, B1 => n4481, B2 => n555
                           , ZN => n5034);
   U3880 : NAND2_X1 port map( A1 => n5036, A2 => n5037, ZN => n5029);
   U3881 : AOI22_X1 port map( A1 => n4484, A2 => n683, B1 => n4485, B2 => n651,
                           ZN => n5037);
   U3882 : AOI22_X1 port map( A1 => n4486, A2 => n715, B1 => n4487, B2 => n587,
                           ZN => n5036);
   U3883 : NAND2_X1 port map( A1 => n5038, A2 => n5039, ZN => n5028);
   U3884 : AOI22_X1 port map( A1 => n5581, A2 => n491, B1 => n5577, B2 => n363,
                           ZN => n5039);
   U3885 : AOI22_X1 port map( A1 => n4492, A2 => n523, B1 => n4493, B2 => n331,
                           ZN => n5038);
   U3886 : NAND2_X1 port map( A1 => n5040, A2 => n5041, ZN => n3175);
   U3887 : NOR4_X1 port map( A1 => n5042, A2 => n5043, A3 => n5044, A4 => n5045
                           , ZN => n5041);
   U3888 : OAI21_X1 port map( B1 => n1445, B2 => n4442, A => n5046, ZN => n5045
                           );
   U3889 : NAND2_X1 port map( A1 => n4444, A2 => n6837, ZN => n5046);
   U3890 : OAI21_X1 port map( B1 => n5523, B2 => n4445, A => n5047, ZN => n5044
                           );
   U3891 : AOI22_X1 port map( A1 => n4447, A2 => n6685, B1 => n4448, B2 => 
                           n6889, ZN => n5047);
   U3892 : NAND2_X1 port map( A1 => n5048, A2 => n5049, ZN => n5043);
   U3893 : AOI22_X1 port map( A1 => n5649, A2 => n2808, B1 => n4452, B2 => 
                           n6888, ZN => n5049);
   U3894 : AOI22_X1 port map( A1 => n4453, A2 => n6626, B1 => n4454, B2 => 
                           n6720, ZN => n5048);
   U3896 : AOI22_X1 port map( A1 => n4459, A2 => n6752, B1 => n4460, B2 => 
                           n6997, ZN => n5053);
   U3897 : AOI22_X1 port map( A1 => n4461, A2 => n6645, B1 => n5629, B2 => 
                           n6887, ZN => n5052);
   U3898 : AOI22_X1 port map( A1 => n4463, A2 => n2175, B1 => n4464, B2 => 
                           n7029, ZN => n5051);
   U3899 : AOI22_X1 port map( A1 => n4465, A2 => n618, B1 => n4466, B2 => n458,
                           ZN => n5050);
   U3900 : NOR4_X1 port map( A1 => n5054, A2 => n5055, A3 => n5056, A4 => n5057
                           , ZN => n5040);
   U3901 : NAND2_X1 port map( A1 => n5058, A2 => n5059, ZN => n5057);
   U3902 : AOI22_X1 port map( A1 => n4473, A2 => n394, B1 => n4474, B2 => n7061
                           , ZN => n5059);
   U3903 : AOI22_X1 port map( A1 => n4475, A2 => n6818, B1 => n5932, B2 => 
                           OUT2_9_port, ZN => n5058);
   U3904 : NAND2_X1 port map( A1 => n5060, A2 => n5061, ZN => n5056);
   U3905 : AOI22_X1 port map( A1 => n5605, A2 => n426, B1 => n5601, B2 => n6961
                           , ZN => n5061);
   U3906 : AOI22_X1 port map( A1 => n4480, A2 => n6786, B1 => n4481, B2 => n554
                           , ZN => n5060);
   U3907 : NAND2_X1 port map( A1 => n5062, A2 => n5063, ZN => n5055);
   U3908 : AOI22_X1 port map( A1 => n4484, A2 => n682, B1 => n4485, B2 => n650,
                           ZN => n5063);
   U3909 : AOI22_X1 port map( A1 => n4486, A2 => n714, B1 => n4487, B2 => n586,
                           ZN => n5062);
   U3910 : NAND2_X1 port map( A1 => n5064, A2 => n5065, ZN => n5054);
   U3911 : AOI22_X1 port map( A1 => n5581, A2 => n490, B1 => n5577, B2 => n362,
                           ZN => n5065);
   U3912 : AOI22_X1 port map( A1 => n4492, A2 => n522, B1 => n4493, B2 => n330,
                           ZN => n5064);
   U3913 : NAND2_X1 port map( A1 => n5066, A2 => n5067, ZN => n3174);
   U3914 : NOR4_X1 port map( A1 => n5068, A2 => n5069, A3 => n5070, A4 => n5071
                           , ZN => n5067);
   U3915 : OAI21_X1 port map( B1 => n1446, B2 => n4442, A => n5072, ZN => n5071
                           );
   U3916 : NAND2_X1 port map( A1 => n4444, A2 => n6836, ZN => n5072);
   U3917 : OAI21_X1 port map( B1 => n6082, B2 => n4445, A => n5073, ZN => n5070
                           );
   U3918 : AOI22_X1 port map( A1 => n4447, A2 => n6684, B1 => n4448, B2 => 
                           n6886, ZN => n5073);
   U3919 : NAND2_X1 port map( A1 => n5074, A2 => n5075, ZN => n5069);
   U3920 : AOI22_X1 port map( A1 => n5649, A2 => n2807, B1 => n4452, B2 => 
                           n6885, ZN => n5075);
   U3921 : AOI22_X1 port map( A1 => n4453, A2 => n6627, B1 => n4454, B2 => 
                           n6719, ZN => n5074);
   U3923 : AOI22_X1 port map( A1 => n4459, A2 => n6751, B1 => n4460, B2 => 
                           n6996, ZN => n5079);
   U3924 : AOI22_X1 port map( A1 => n4461, A2 => n6644, B1 => n5629, B2 => 
                           n6884, ZN => n5078);
   U3925 : AOI22_X1 port map( A1 => n4463, A2 => n2170, B1 => n4464, B2 => 
                           n7028, ZN => n5077);
   U3926 : AOI22_X1 port map( A1 => n4465, A2 => n617, B1 => n4466, B2 => n457,
                           ZN => n5076);
   U3927 : NOR4_X1 port map( A1 => n5080, A2 => n5081, A3 => n5082, A4 => n5083
                           , ZN => n5066);
   U3928 : NAND2_X1 port map( A1 => n5084, A2 => n5085, ZN => n5083);
   U3929 : AOI22_X1 port map( A1 => n4473, A2 => n393, B1 => n4474, B2 => n7060
                           , ZN => n5085);
   U3930 : AOI22_X1 port map( A1 => n4475, A2 => n6819, B1 => n5934, B2 => 
                           OUT2_8_port, ZN => n5084);
   U3931 : NAND2_X1 port map( A1 => n5086, A2 => n5087, ZN => n5082);
   U3932 : AOI22_X1 port map( A1 => n5605, A2 => n425, B1 => n5601, B2 => n6962
                           , ZN => n5087);
   U3933 : AOI22_X1 port map( A1 => n4480, A2 => n6787, B1 => n4481, B2 => n553
                           , ZN => n5086);
   U3934 : NAND2_X1 port map( A1 => n5088, A2 => n5089, ZN => n5081);
   U3935 : AOI22_X1 port map( A1 => n4484, A2 => n681, B1 => n4485, B2 => n649,
                           ZN => n5089);
   U3936 : AOI22_X1 port map( A1 => n4486, A2 => n713, B1 => n4487, B2 => n585,
                           ZN => n5088);
   U3937 : NAND2_X1 port map( A1 => n5090, A2 => n5091, ZN => n5080);
   U3938 : AOI22_X1 port map( A1 => n5581, A2 => n489, B1 => n5577, B2 => n361,
                           ZN => n5091);
   U3939 : AOI22_X1 port map( A1 => n4492, A2 => n521, B1 => n4493, B2 => n329,
                           ZN => n5090);
   U3940 : NAND2_X1 port map( A1 => n5092, A2 => n5093, ZN => n3173);
   U3941 : NOR4_X1 port map( A1 => n5094, A2 => n5095, A3 => n5096, A4 => n5097
                           , ZN => n5093);
   U3942 : OAI21_X1 port map( B1 => n1447, B2 => n4442, A => n5098, ZN => n5097
                           );
   U3943 : NAND2_X1 port map( A1 => n4444, A2 => n6835, ZN => n5098);
   U3944 : OAI21_X1 port map( B1 => n6083, B2 => n4445, A => n5099, ZN => n5096
                           );
   U3945 : AOI22_X1 port map( A1 => n4447, A2 => n6683, B1 => n4448, B2 => 
                           n6883, ZN => n5099);
   U3946 : NAND2_X1 port map( A1 => n5100, A2 => n5101, ZN => n5095);
   U3947 : AOI22_X1 port map( A1 => n5649, A2 => n6675, B1 => n4452, B2 => 
                           n6882, ZN => n5101);
   U3948 : AOI22_X1 port map( A1 => n4453, A2 => n6628, B1 => n4454, B2 => 
                           n6718, ZN => n5100);
   U3950 : AOI22_X1 port map( A1 => n4459, A2 => n6750, B1 => n4460, B2 => 
                           n6995, ZN => n5105);
   U3951 : AOI22_X1 port map( A1 => n4461, A2 => n6643, B1 => n5629, B2 => 
                           n6881, ZN => n5104);
   U3952 : AOI22_X1 port map( A1 => n4463, A2 => n2165, B1 => n4464, B2 => 
                           n7027, ZN => n5103);
   U3953 : AOI22_X1 port map( A1 => n4465, A2 => n616, B1 => n4466, B2 => n456,
                           ZN => n5102);
   U3954 : NOR4_X1 port map( A1 => n5106, A2 => n5107, A3 => n5108, A4 => n5109
                           , ZN => n5092);
   U3955 : NAND2_X1 port map( A1 => n5110, A2 => n5111, ZN => n5109);
   U3956 : AOI22_X1 port map( A1 => n4473, A2 => n392, B1 => n4474, B2 => n7059
                           , ZN => n5111);
   U3957 : AOI22_X1 port map( A1 => n4475, A2 => n6820, B1 => n5935, B2 => 
                           OUT2_7_port, ZN => n5110);
   U3958 : NAND2_X1 port map( A1 => n5112, A2 => n5113, ZN => n5108);
   U3959 : AOI22_X1 port map( A1 => n5605, A2 => n424, B1 => n5601, B2 => n6963
                           , ZN => n5113);
   U3960 : AOI22_X1 port map( A1 => n4480, A2 => n6788, B1 => n4481, B2 => n552
                           , ZN => n5112);
   U3961 : NAND2_X1 port map( A1 => n5114, A2 => n5115, ZN => n5107);
   U3962 : AOI22_X1 port map( A1 => n4484, A2 => n680, B1 => n4485, B2 => n648,
                           ZN => n5115);
   U3963 : AOI22_X1 port map( A1 => n4486, A2 => n712, B1 => n4487, B2 => n584,
                           ZN => n5114);
   U3964 : NAND2_X1 port map( A1 => n5116, A2 => n5117, ZN => n5106);
   U3965 : AOI22_X1 port map( A1 => n5581, A2 => n488, B1 => n5577, B2 => n360,
                           ZN => n5117);
   U3966 : AOI22_X1 port map( A1 => n4492, A2 => n520, B1 => n4493, B2 => n328,
                           ZN => n5116);
   U3967 : NAND2_X1 port map( A1 => n5118, A2 => n5119, ZN => n3172);
   U3968 : NOR4_X1 port map( A1 => n5120, A2 => n5121, A3 => n5122, A4 => n5123
                           , ZN => n5119);
   U3969 : OAI21_X1 port map( B1 => n1448, B2 => n4442, A => n5124, ZN => n5123
                           );
   U3970 : NAND2_X1 port map( A1 => n4444, A2 => n6834, ZN => n5124);
   U3971 : OAI21_X1 port map( B1 => n6084, B2 => n4445, A => n5125, ZN => n5122
                           );
   U3972 : AOI22_X1 port map( A1 => n4447, A2 => n6682, B1 => n4448, B2 => 
                           n6880, ZN => n5125);
   U3973 : NAND2_X1 port map( A1 => n5126, A2 => n5127, ZN => n5121);
   U3974 : AOI22_X1 port map( A1 => n5649, A2 => n6674, B1 => n4452, B2 => 
                           n6879, ZN => n5127);
   U3975 : AOI22_X1 port map( A1 => n4453, A2 => n6629, B1 => n4454, B2 => 
                           n6717, ZN => n5126);
   U3977 : AOI22_X1 port map( A1 => n4459, A2 => n6749, B1 => n4460, B2 => 
                           n6994, ZN => n5131);
   U3978 : AOI22_X1 port map( A1 => n4461, A2 => n6642, B1 => n5629, B2 => 
                           n6878, ZN => n5130);
   U3979 : AOI22_X1 port map( A1 => n4463, A2 => n2160, B1 => n4464, B2 => 
                           n7026, ZN => n5129);
   U3980 : AOI22_X1 port map( A1 => n4465, A2 => n615, B1 => n4466, B2 => n455,
                           ZN => n5128);
   U3981 : NOR4_X1 port map( A1 => n5132, A2 => n5133, A3 => n5134, A4 => n5135
                           , ZN => n5118);
   U3982 : NAND2_X1 port map( A1 => n5136, A2 => n5137, ZN => n5135);
   U3983 : AOI22_X1 port map( A1 => n4473, A2 => n391, B1 => n4474, B2 => n7058
                           , ZN => n5137);
   U3984 : AOI22_X1 port map( A1 => n4475, A2 => n6821, B1 => n5934, B2 => 
                           OUT2_6_port, ZN => n5136);
   U3985 : NAND2_X1 port map( A1 => n5138, A2 => n5139, ZN => n5134);
   U3986 : AOI22_X1 port map( A1 => n5605, A2 => n423, B1 => n5601, B2 => n6964
                           , ZN => n5139);
   U3987 : AOI22_X1 port map( A1 => n4480, A2 => n6789, B1 => n4481, B2 => n551
                           , ZN => n5138);
   U3988 : NAND2_X1 port map( A1 => n5140, A2 => n5141, ZN => n5133);
   U3989 : AOI22_X1 port map( A1 => n4484, A2 => n679, B1 => n4485, B2 => n647,
                           ZN => n5141);
   U3990 : AOI22_X1 port map( A1 => n4486, A2 => n711, B1 => n4487, B2 => n583,
                           ZN => n5140);
   U3991 : NAND2_X1 port map( A1 => n5142, A2 => n5143, ZN => n5132);
   U3992 : AOI22_X1 port map( A1 => n5581, A2 => n487, B1 => n5577, B2 => n359,
                           ZN => n5143);
   U3993 : AOI22_X1 port map( A1 => n4492, A2 => n519, B1 => n4493, B2 => n327,
                           ZN => n5142);
   U3994 : NAND2_X1 port map( A1 => n5144, A2 => n5145, ZN => n3171);
   U3995 : NOR4_X1 port map( A1 => n5146, A2 => n5147, A3 => n5148, A4 => n5149
                           , ZN => n5145);
   U3996 : OAI21_X1 port map( B1 => n1449, B2 => n4442, A => n5150, ZN => n5149
                           );
   U3997 : NAND2_X1 port map( A1 => n5663, A2 => n6833, ZN => n5150);
   U3998 : OAI21_X1 port map( B1 => n6085, B2 => n4445, A => n5151, ZN => n5148
                           );
   U3999 : AOI22_X1 port map( A1 => n5657, A2 => n6681, B1 => n5654, B2 => 
                           n6877, ZN => n5151);
   U4000 : NAND2_X1 port map( A1 => n5152, A2 => n5153, ZN => n5147);
   U4001 : AOI22_X1 port map( A1 => n5649, A2 => n6673, B1 => n4452, B2 => 
                           n6876, ZN => n5153);
   U4002 : AOI22_X1 port map( A1 => n5645, A2 => n6630, B1 => n5642, B2 => 
                           n6716, ZN => n5152);
   U4004 : AOI22_X1 port map( A1 => n5639, A2 => n6748, B1 => n4460, B2 => 
                           n6993, ZN => n5157);
   U4005 : AOI22_X1 port map( A1 => n5633, A2 => n6641, B1 => n4462, B2 => 
                           n6875, ZN => n5156);
   U4006 : AOI22_X1 port map( A1 => n5627, A2 => n2155, B1 => n4464, B2 => 
                           n7025, ZN => n5155);
   U4007 : AOI22_X1 port map( A1 => n5621, A2 => n614, B1 => n5618, B2 => n454,
                           ZN => n5154);
   U4008 : NOR4_X1 port map( A1 => n5158, A2 => n5159, A3 => n5160, A4 => n5161
                           , ZN => n5144);
   U4009 : NAND2_X1 port map( A1 => n5162, A2 => n5163, ZN => n5161);
   U4010 : AOI22_X1 port map( A1 => n5615, A2 => n390, B1 => n5612, B2 => n7057
                           , ZN => n5163);
   U4011 : AOI22_X1 port map( A1 => n5609, A2 => n6822, B1 => n5935, B2 => 
                           OUT2_5_port, ZN => n5162);
   U4012 : NAND2_X1 port map( A1 => n5164, A2 => n5165, ZN => n5160);
   U4013 : AOI22_X1 port map( A1 => n5605, A2 => n422, B1 => n5601, B2 => n6965
                           , ZN => n5165);
   U4014 : AOI22_X1 port map( A1 => n5600, A2 => n6790, B1 => n5597, B2 => n550
                           , ZN => n5164);
   U4015 : NAND2_X1 port map( A1 => n5166, A2 => n5167, ZN => n5159);
   U4016 : AOI22_X1 port map( A1 => n4484, A2 => n678, B1 => n5591, B2 => n646,
                           ZN => n5167);
   U4017 : AOI22_X1 port map( A1 => n5588, A2 => n710, B1 => n5585, B2 => n582,
                           ZN => n5166);
   U4018 : NAND2_X1 port map( A1 => n5168, A2 => n5169, ZN => n5158);
   U4019 : AOI22_X1 port map( A1 => n5581, A2 => n486, B1 => n5577, B2 => n358,
                           ZN => n5169);
   U4020 : AOI22_X1 port map( A1 => n5576, A2 => n518, B1 => n5573, B2 => n326,
                           ZN => n5168);
   U4021 : NAND2_X1 port map( A1 => n5170, A2 => n5171, ZN => n3170);
   U4022 : NOR4_X1 port map( A1 => n5172, A2 => n5173, A3 => n5174, A4 => n5175
                           , ZN => n5171);
   U4023 : OAI21_X1 port map( B1 => n1450, B2 => n4442, A => n5176, ZN => n5175
                           );
   U4024 : NAND2_X1 port map( A1 => n5663, A2 => n6832, ZN => n5176);
   U4025 : OAI21_X1 port map( B1 => n6086, B2 => n4445, A => n5177, ZN => n5174
                           );
   U4026 : AOI22_X1 port map( A1 => n5657, A2 => n6680, B1 => n5654, B2 => 
                           n6874, ZN => n5177);
   U4027 : NAND2_X1 port map( A1 => n5178, A2 => n5179, ZN => n5173);
   U4028 : AOI22_X1 port map( A1 => n5649, A2 => n6672, B1 => n5648, B2 => 
                           n6873, ZN => n5179);
   U4029 : AOI22_X1 port map( A1 => n5645, A2 => n6631, B1 => n5642, B2 => 
                           n6715, ZN => n5178);
   U4031 : AOI22_X1 port map( A1 => n5639, A2 => n6747, B1 => n5636, B2 => 
                           n6992, ZN => n5183);
   U4032 : AOI22_X1 port map( A1 => n5633, A2 => n6640, B1 => n4462, B2 => 
                           n6872, ZN => n5182);
   U4033 : AOI22_X1 port map( A1 => n5627, A2 => n2150, B1 => n5624, B2 => 
                           n7024, ZN => n5181);
   U4034 : AOI22_X1 port map( A1 => n5621, A2 => n613, B1 => n5618, B2 => n453,
                           ZN => n5180);
   U4035 : NOR4_X1 port map( A1 => n5184, A2 => n5185, A3 => n5186, A4 => n5187
                           , ZN => n5170);
   U4036 : NAND2_X1 port map( A1 => n5188, A2 => n5189, ZN => n5187);
   U4037 : AOI22_X1 port map( A1 => n5615, A2 => n389, B1 => n5612, B2 => n7056
                           , ZN => n5189);
   U4038 : AOI22_X1 port map( A1 => n5609, A2 => n6823, B1 => n5934, B2 => 
                           OUT2_4_port, ZN => n5188);
   U4039 : NAND2_X1 port map( A1 => n5190, A2 => n5191, ZN => n5186);
   U4040 : AOI22_X1 port map( A1 => n4478, A2 => n421, B1 => n5601, B2 => n6966
                           , ZN => n5191);
   U4041 : AOI22_X1 port map( A1 => n5600, A2 => n6791, B1 => n5597, B2 => n549
                           , ZN => n5190);
   U4042 : NAND2_X1 port map( A1 => n5192, A2 => n5193, ZN => n5185);
   U4043 : AOI22_X1 port map( A1 => n5594, A2 => n677, B1 => n5591, B2 => n645,
                           ZN => n5193);
   U4044 : AOI22_X1 port map( A1 => n5588, A2 => n709, B1 => n5585, B2 => n581,
                           ZN => n5192);
   U4045 : NAND2_X1 port map( A1 => n5194, A2 => n5195, ZN => n5184);
   U4046 : AOI22_X1 port map( A1 => n4490, A2 => n485, B1 => n5577, B2 => n357,
                           ZN => n5195);
   U4047 : AOI22_X1 port map( A1 => n5576, A2 => n517, B1 => n5573, B2 => n325,
                           ZN => n5194);
   U4048 : NAND2_X1 port map( A1 => n5196, A2 => n5197, ZN => n3169);
   U4049 : NOR4_X1 port map( A1 => n5198, A2 => n5199, A3 => n5200, A4 => n5201
                           , ZN => n5197);
   U4050 : OAI21_X1 port map( B1 => n1451, B2 => n5666, A => n5202, ZN => n5201
                           );
   U4051 : NAND2_X1 port map( A1 => n5663, A2 => n6831, ZN => n5202);
   U4052 : OAI21_X1 port map( B1 => n6087, B2 => n5660, A => n5203, ZN => n5200
                           );
   U4053 : AOI22_X1 port map( A1 => n5657, A2 => n6679, B1 => n5654, B2 => 
                           n6871, ZN => n5203);
   U4054 : NAND2_X1 port map( A1 => n5204, A2 => n5205, ZN => n5199);
   U4055 : AOI22_X1 port map( A1 => n5649, A2 => n6671, B1 => n5648, B2 => 
                           n6870, ZN => n5205);
   U4056 : AOI22_X1 port map( A1 => n5645, A2 => n6632, B1 => n5642, B2 => 
                           n6714, ZN => n5204);
   U4058 : AOI22_X1 port map( A1 => n5639, A2 => n6746, B1 => n5636, B2 => 
                           n6991, ZN => n5209);
   U4059 : AOI22_X1 port map( A1 => n5633, A2 => n6639, B1 => n4462, B2 => 
                           n6869, ZN => n5208);
   U4060 : AOI22_X1 port map( A1 => n5627, A2 => n2145, B1 => n5624, B2 => 
                           n7023, ZN => n5207);
   U4061 : AOI22_X1 port map( A1 => n5621, A2 => n612, B1 => n5618, B2 => n452,
                           ZN => n5206);
   U4062 : NOR4_X1 port map( A1 => n5210, A2 => n5211, A3 => n5212, A4 => n5213
                           , ZN => n5196);
   U4063 : NAND2_X1 port map( A1 => n5214, A2 => n5215, ZN => n5213);
   U4064 : AOI22_X1 port map( A1 => n5615, A2 => n388, B1 => n5612, B2 => n7055
                           , ZN => n5215);
   U4065 : AOI22_X1 port map( A1 => n5609, A2 => n6824, B1 => n5932, B2 => 
                           OUT2_3_port, ZN => n5214);
   U4066 : NAND2_X1 port map( A1 => n5216, A2 => n5217, ZN => n5212);
   U4067 : AOI22_X1 port map( A1 => n4478, A2 => n420, B1 => n5601, B2 => n6967
                           , ZN => n5217);
   U4068 : AOI22_X1 port map( A1 => n5600, A2 => n6792, B1 => n5597, B2 => n548
                           , ZN => n5216);
   U4069 : NAND2_X1 port map( A1 => n5218, A2 => n5219, ZN => n5211);
   U4070 : AOI22_X1 port map( A1 => n5594, A2 => n676, B1 => n5591, B2 => n644,
                           ZN => n5219);
   U4071 : AOI22_X1 port map( A1 => n5588, A2 => n708, B1 => n5585, B2 => n580,
                           ZN => n5218);
   U4072 : NAND2_X1 port map( A1 => n5220, A2 => n5221, ZN => n5210);
   U4073 : AOI22_X1 port map( A1 => n4490, A2 => n484, B1 => n5577, B2 => n356,
                           ZN => n5221);
   U4074 : AOI22_X1 port map( A1 => n5576, A2 => n516, B1 => n5573, B2 => n324,
                           ZN => n5220);
   U4075 : NAND2_X1 port map( A1 => n5222, A2 => n5223, ZN => n3168);
   U4076 : NOR4_X1 port map( A1 => n5224, A2 => n5225, A3 => n5226, A4 => n5227
                           , ZN => n5223);
   U4077 : OAI21_X1 port map( B1 => n1452, B2 => n5666, A => n5228, ZN => n5227
                           );
   U4078 : NAND2_X1 port map( A1 => n5663, A2 => n6830, ZN => n5228);
   U4079 : OAI21_X1 port map( B1 => n6088, B2 => n5660, A => n5229, ZN => n5226
                           );
   U4080 : AOI22_X1 port map( A1 => n5657, A2 => n6678, B1 => n5654, B2 => 
                           n6868, ZN => n5229);
   U4081 : NAND2_X1 port map( A1 => n5230, A2 => n5231, ZN => n5225);
   U4082 : AOI22_X1 port map( A1 => n5649, A2 => n6670, B1 => n5648, B2 => 
                           n6867, ZN => n5231);
   U4083 : AOI22_X1 port map( A1 => n5645, A2 => n6633, B1 => n5642, B2 => 
                           n6713, ZN => n5230);
   U4085 : AOI22_X1 port map( A1 => n5639, A2 => n6745, B1 => n5636, B2 => 
                           n6990, ZN => n5235);
   U4086 : AOI22_X1 port map( A1 => n5633, A2 => n6638, B1 => n4462, B2 => 
                           n6866, ZN => n5234);
   U4087 : AOI22_X1 port map( A1 => n5627, A2 => n2140, B1 => n5624, B2 => 
                           n7022, ZN => n5233);
   U4088 : AOI22_X1 port map( A1 => n5621, A2 => n611, B1 => n5618, B2 => n451,
                           ZN => n5232);
   U4089 : NOR4_X1 port map( A1 => n5236, A2 => n5237, A3 => n5238, A4 => n5239
                           , ZN => n5222);
   U4090 : NAND2_X1 port map( A1 => n5240, A2 => n5241, ZN => n5239);
   U4091 : AOI22_X1 port map( A1 => n5615, A2 => n387, B1 => n5612, B2 => n7054
                           , ZN => n5241);
   U4092 : AOI22_X1 port map( A1 => n5609, A2 => n6825, B1 => n5935, B2 => 
                           OUT2_2_port, ZN => n5240);
   U4093 : NAND2_X1 port map( A1 => n5242, A2 => n5243, ZN => n5238);
   U4094 : AOI22_X1 port map( A1 => n4478, A2 => n419, B1 => n5601, B2 => n6968
                           , ZN => n5243);
   U4095 : AOI22_X1 port map( A1 => n5600, A2 => n6793, B1 => n5597, B2 => n547
                           , ZN => n5242);
   U4096 : NAND2_X1 port map( A1 => n5244, A2 => n5245, ZN => n5237);
   U4097 : AOI22_X1 port map( A1 => n5594, A2 => n675, B1 => n5591, B2 => n643,
                           ZN => n5245);
   U4098 : AOI22_X1 port map( A1 => n5588, A2 => n707, B1 => n5585, B2 => n579,
                           ZN => n5244);
   U4099 : NAND2_X1 port map( A1 => n5246, A2 => n5247, ZN => n5236);
   U4100 : AOI22_X1 port map( A1 => n4490, A2 => n483, B1 => n5577, B2 => n355,
                           ZN => n5247);
   U4101 : AOI22_X1 port map( A1 => n5576, A2 => n515, B1 => n5573, B2 => n323,
                           ZN => n5246);
   U4102 : NAND2_X1 port map( A1 => n5248, A2 => n5249, ZN => n3167);
   U4103 : NOR4_X1 port map( A1 => n5250, A2 => n5251, A3 => n5252, A4 => n5253
                           , ZN => n5249);
   U4104 : OAI21_X1 port map( B1 => n1453, B2 => n5666, A => n5254, ZN => n5253
                           );
   U4105 : NAND2_X1 port map( A1 => n5663, A2 => n6829, ZN => n5254);
   U4106 : OAI21_X1 port map( B1 => n6089, B2 => n5660, A => n5255, ZN => n5252
                           );
   U4107 : AOI22_X1 port map( A1 => n5657, A2 => n6677, B1 => n5654, B2 => 
                           n6865, ZN => n5255);
   U4108 : NAND2_X1 port map( A1 => n5256, A2 => n5257, ZN => n5251);
   U4109 : AOI22_X1 port map( A1 => n5649, A2 => n6669, B1 => n5648, B2 => 
                           n6864, ZN => n5257);
   U4110 : AOI22_X1 port map( A1 => n5645, A2 => n6634, B1 => n5642, B2 => 
                           n6712, ZN => n5256);
   U4112 : AOI22_X1 port map( A1 => n5639, A2 => n6744, B1 => n5636, B2 => 
                           n6989, ZN => n5261);
   U4113 : AOI22_X1 port map( A1 => n5633, A2 => n6637, B1 => n4462, B2 => 
                           n6863, ZN => n5260);
   U4114 : AOI22_X1 port map( A1 => n5627, A2 => n2135, B1 => n5624, B2 => 
                           n7021, ZN => n5259);
   U4115 : AOI22_X1 port map( A1 => n5621, A2 => n610, B1 => n5618, B2 => n450,
                           ZN => n5258);
   U4116 : NOR4_X1 port map( A1 => n5262, A2 => n5263, A3 => n5264, A4 => n5265
                           , ZN => n5248);
   U4117 : NAND2_X1 port map( A1 => n5266, A2 => n5267, ZN => n5265);
   U4118 : AOI22_X1 port map( A1 => n5615, A2 => n386, B1 => n5612, B2 => n7053
                           , ZN => n5267);
   U4119 : AOI22_X1 port map( A1 => n5609, A2 => n6826, B1 => n5934, B2 => 
                           OUT2_1_port, ZN => n5266);
   U4120 : NAND2_X1 port map( A1 => n5268, A2 => n5269, ZN => n5264);
   U4121 : AOI22_X1 port map( A1 => n4478, A2 => n418, B1 => n5601, B2 => n6969
                           , ZN => n5269);
   U4122 : AOI22_X1 port map( A1 => n5600, A2 => n6794, B1 => n5597, B2 => n546
                           , ZN => n5268);
   U4123 : NAND2_X1 port map( A1 => n5270, A2 => n5271, ZN => n5263);
   U4124 : AOI22_X1 port map( A1 => n5594, A2 => n674, B1 => n5591, B2 => n642,
                           ZN => n5271);
   U4125 : AOI22_X1 port map( A1 => n5588, A2 => n706, B1 => n5585, B2 => n578,
                           ZN => n5270);
   U4126 : NAND2_X1 port map( A1 => n5272, A2 => n5273, ZN => n5262);
   U4127 : AOI22_X1 port map( A1 => n4490, A2 => n482, B1 => n5577, B2 => n354,
                           ZN => n5273);
   U4128 : AOI22_X1 port map( A1 => n5576, A2 => n514, B1 => n5573, B2 => n322,
                           ZN => n5272);
   U4129 : NAND2_X1 port map( A1 => n5274, A2 => n5275, ZN => n3166);
   U4130 : NOR4_X1 port map( A1 => n5276, A2 => n5277, A3 => n5278, A4 => n5279
                           , ZN => n5275);
   U4131 : OAI21_X1 port map( B1 => n1454, B2 => n5666, A => n5280, ZN => n5279
                           );
   U4132 : NAND2_X1 port map( A1 => n5663, A2 => n6828, ZN => n5280);
   U4133 : NOR2_X1 port map( A1 => n5281, A2 => n5282, ZN => n4444);
   U4134 : OR2_X1 port map( A1 => n5281, A2 => n5283, ZN => n4442);
   U4135 : OAI21_X1 port map( B1 => n6090, B2 => n5660, A => n5284, ZN => n5278
                           );
   U4136 : AOI22_X1 port map( A1 => n5657, A2 => n6676, B1 => n5654, B2 => 
                           n6862, ZN => n5284);
   U4137 : NOR2_X1 port map( A1 => n5283, A2 => n5285, ZN => n4448);
   U4138 : NOR2_X1 port map( A1 => n5285, A2 => n5282, ZN => n4447);
   U4139 : NAND2_X1 port map( A1 => n5286, A2 => n5287, ZN => n4445);
   U4140 : NOR4_X1 port map( A1 => n6603, A2 => n5288, A3 => n5289, A4 => n5290
                           , ZN => n5287);
   U4141 : NOR3_X1 port map( A1 => n5291, A2 => n5292, A3 => n5293, ZN => n5286
                           );
   U4142 : NAND2_X1 port map( A1 => n5294, A2 => n5295, ZN => n5277);
   U4143 : AOI22_X1 port map( A1 => n5649, A2 => n6668, B1 => n5648, B2 => 
                           n6861, ZN => n5295);
   U4144 : NOR2_X1 port map( A1 => n5296, A2 => n5297, ZN => n4452);
   U4145 : NOR2_X1 port map( A1 => n5297, A2 => n5298, ZN => n4451);
   U4146 : AOI22_X1 port map( A1 => n5645, A2 => n6635, B1 => n5642, B2 => 
                           n6711, ZN => n5294);
   U4147 : NOR2_X1 port map( A1 => n5299, A2 => n5296, ZN => n4454);
   U4148 : NOR2_X1 port map( A1 => n5297, A2 => n5283, ZN => n4453);
   U4150 : AOI22_X1 port map( A1 => n5639, A2 => n6743, B1 => n5636, B2 => 
                           n6988, ZN => n5303);
   U4151 : NOR2_X1 port map( A1 => n5304, A2 => n5281, ZN => n4460);
   U4152 : NOR2_X1 port map( A1 => n5305, A2 => n5281, ZN => n4459);
   U4153 : AOI22_X1 port map( A1 => n5633, A2 => n6636, B1 => n5629, B2 => 
                           n6860, ZN => n5302);
   U4154 : NOR2_X1 port map( A1 => n5299, A2 => n5298, ZN => n4462);
   U4155 : NOR2_X1 port map( A1 => n5299, A2 => n5306, ZN => n4461);
   U4156 : AOI22_X1 port map( A1 => n5627, A2 => n2130, B1 => n5624, B2 => 
                           n7020, ZN => n5301);
   U4157 : NOR2_X1 port map( A1 => n5305, A2 => n5285, ZN => n4464);
   U4158 : NOR2_X1 port map( A1 => n5304, A2 => n5285, ZN => n4463);
   U4159 : AOI22_X1 port map( A1 => n5621, A2 => n609, B1 => n5618, B2 => n449,
                           ZN => n5300);
   U4160 : NOR2_X1 port map( A1 => n5307, A2 => n5281, ZN => n4466);
   U4161 : NOR2_X1 port map( A1 => n5307, A2 => n5297, ZN => n4465);
   U4162 : NOR4_X1 port map( A1 => n5308, A2 => n5309, A3 => n5310, A4 => n5311
                           , ZN => n5274);
   U4163 : NAND2_X1 port map( A1 => n5312, A2 => n5313, ZN => n5311);
   U4164 : AOI22_X1 port map( A1 => n5615, A2 => n385, B1 => n5612, B2 => n7052
                           , ZN => n5313);
   U4165 : NOR2_X1 port map( A1 => n5307, A2 => n5299, ZN => n4474);
   U4166 : NOR2_X1 port map( A1 => n5304, A2 => n5299, ZN => n4473);
   U4167 : AOI22_X1 port map( A1 => n5609, A2 => n6827, B1 => n5935, B2 => 
                           OUT2_0_port, ZN => n5312);
   U4168 : NOR2_X1 port map( A1 => n5305, A2 => n5299, ZN => n4475);
   U4169 : NAND2_X1 port map( A1 => n5314, A2 => n5315, ZN => n5310);
   U4170 : AOI22_X1 port map( A1 => n4478, A2 => n417, B1 => n5601, B2 => n6970
                           , ZN => n5315);
   U4171 : NOR2_X1 port map( A1 => n5285, A2 => n5306, ZN => n4479);
   U4172 : NOR2_X1 port map( A1 => n5305, A2 => n5297, ZN => n4478);
   U4173 : NAND2_X1 port map( A1 => n5316, A2 => ADD_RD2(3), ZN => n5305);
   U4174 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => n6058, ZN => n5316);
   U4175 : AOI22_X1 port map( A1 => n5600, A2 => n6795, B1 => n5597, B2 => n545
                           , ZN => n5314);
   U4176 : NOR2_X1 port map( A1 => n5304, A2 => n5297, ZN => n4481);
   U4177 : NAND2_X1 port map( A1 => n5317, A2 => ADD_RD2(3), ZN => n5304);
   U4178 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(0), ZN => n5317);
   U4179 : NOR2_X1 port map( A1 => n5281, A2 => n5306, ZN => n4480);
   U4180 : NAND2_X1 port map( A1 => n5318, A2 => n5319, ZN => n5309);
   U4181 : AOI22_X1 port map( A1 => n5594, A2 => n673, B1 => n5591, B2 => n641,
                           ZN => n5319);
   U4182 : NOR2_X1 port map( A1 => n5298, A2 => n5285, ZN => n4485);
   U4183 : NOR2_X1 port map( A1 => n5297, A2 => n5282, ZN => n4484);
   U4184 : NAND2_X1 port map( A1 => n5320, A2 => n5321, ZN => n5297);
   U4185 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), ZN => n5320);
   U4186 : AOI22_X1 port map( A1 => n5588, A2 => n705, B1 => n5585, B2 => n577,
                           ZN => n5318);
   U4187 : NOR2_X1 port map( A1 => n5307, A2 => n5285, ZN => n4487);
   U4188 : OR2_X1 port map( A1 => n5322, A2 => n6058, ZN => n5307);
   U4189 : OR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n5322);
   U4190 : NOR2_X1 port map( A1 => n5299, A2 => n5282, ZN => n4486);
   U4191 : OR2_X1 port map( A1 => n5323, A2 => n6055, ZN => n5282);
   U4192 : OR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(0), ZN => n5323);
   U4193 : NAND2_X1 port map( A1 => n5324, A2 => n5325, ZN => n5308);
   U4194 : AOI22_X1 port map( A1 => n4490, A2 => n481, B1 => n5577, B2 => n353,
                           ZN => n5325);
   U4195 : NOR2_X1 port map( A1 => n5296, A2 => n5281, ZN => n4491);
   U4196 : NOR2_X1 port map( A1 => n5296, A2 => n5285, ZN => n4490);
   U4197 : NAND2_X1 port map( A1 => n5326, A2 => n5321, ZN => n5285);
   U4198 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => n6057, ZN => n5326);
   U4199 : NAND2_X1 port map( A1 => n5327, A2 => ADD_RD2(3), ZN => n5296);
   U4200 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => n6055, ZN => n5327);
   U4201 : AOI22_X1 port map( A1 => n5576, A2 => n513, B1 => n5573, B2 => n321,
                           ZN => n5324);
   U4202 : NOR2_X1 port map( A1 => n5298, A2 => n5281, ZN => n4493);
   U4203 : NAND2_X1 port map( A1 => n5328, A2 => n5321, ZN => n5281);
   U4204 : NOR2_X1 port map( A1 => n6056, A2 => n6057, ZN => n5328);
   U4205 : NAND2_X1 port map( A1 => n5329, A2 => ADD_RD2(3), ZN => n5298);
   U4206 : NOR2_X1 port map( A1 => n6055, A2 => n6058, ZN => n5329);
   U4207 : NOR2_X1 port map( A1 => n5299, A2 => n5283, ZN => n4492);
   U4208 : OR2_X1 port map( A1 => n5330, A2 => n6058, ZN => n5283);
   U4209 : OR2_X1 port map( A1 => ADD_RD2(3), A2 => n6055, ZN => n5330);
   U4210 : NAND2_X1 port map( A1 => n5331, A2 => n5321, ZN => n5299);
   U4211 : NOR2_X1 port map( A1 => n5291, A2 => n5332, ZN => n5321);
   U4214 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD2(3), Z => n5288);
   U4215 : XOR2_X1 port map( A => ADD_RD2(1), B => ADD_WR(1), Z => n5289);
   U4217 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD2(4), Z => n5292);
   U4218 : XOR2_X1 port map( A => ADD_RD2(0), B => ADD_WR(0), Z => n5290);
   U4219 : XOR2_X1 port map( A => ADD_RD2(2), B => ADD_WR(2), Z => n5293);
   U4220 : NAND2_X1 port map( A1 => n5335, A2 => RD2, ZN => n5291);
   U4221 : NOR2_X1 port map( A1 => n5336, A2 => n5932, ZN => n5335);
   U4222 : NOR3_X1 port map( A1 => n5306, A2 => ADD_RD2(2), A3 => ADD_RD2(1), 
                           ZN => n5336);
   U4223 : NAND2_X1 port map( A1 => n5337, A2 => n6058, ZN => n5306);
   U4224 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n5337);
   U4225 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => n6056, ZN => n5331);
   U4226 : OAI21_X1 port map( B1 => n6076, B2 => n5869, A => n5338, ZN => n3165
                           );
   U4227 : NAND2_X1 port map( A1 => n1828, A2 => n6904, ZN => n5338);
   U4228 : OAI21_X1 port map( B1 => n6077, B2 => n5869, A => n5339, ZN => n3164
                           );
   U4229 : NAND2_X1 port map( A1 => n1828, A2 => n6901, ZN => n5339);
   U4230 : OAI21_X1 port map( B1 => n6078, B2 => n5869, A => n5340, ZN => n3163
                           );
   U4231 : NAND2_X1 port map( A1 => n1828, A2 => n6898, ZN => n5340);
   U4232 : OAI21_X1 port map( B1 => n6079, B2 => n5869, A => n5341, ZN => n3162
                           );
   U4233 : NAND2_X1 port map( A1 => n1828, A2 => n6895, ZN => n5341);
   U4234 : OAI21_X1 port map( B1 => n6080, B2 => n5869, A => n5342, ZN => n3161
                           );
   U4235 : NAND2_X1 port map( A1 => n1828, A2 => n6892, ZN => n5342);
   U4236 : OAI21_X1 port map( B1 => n5523, B2 => n5869, A => n5343, ZN => n3160
                           );
   U4237 : NAND2_X1 port map( A1 => n1828, A2 => n6889, ZN => n5343);
   U4238 : OAI21_X1 port map( B1 => n6082, B2 => n5869, A => n5344, ZN => n3159
                           );
   U4239 : NAND2_X1 port map( A1 => n1828, A2 => n6886, ZN => n5344);
   U4240 : OAI21_X1 port map( B1 => n6083, B2 => n5869, A => n5345, ZN => n3158
                           );
   U4241 : NAND2_X1 port map( A1 => n1828, A2 => n6883, ZN => n5345);
   U4242 : OAI21_X1 port map( B1 => n6084, B2 => n5869, A => n5346, ZN => n3157
                           );
   U4243 : NAND2_X1 port map( A1 => n1828, A2 => n6880, ZN => n5346);
   U4244 : OAI21_X1 port map( B1 => n6085, B2 => n5869, A => n5347, ZN => n3156
                           );
   U4245 : NAND2_X1 port map( A1 => n1828, A2 => n6877, ZN => n5347);
   U4246 : OAI21_X1 port map( B1 => n6086, B2 => n5869, A => n5348, ZN => n3155
                           );
   U4247 : NAND2_X1 port map( A1 => n1828, A2 => n6874, ZN => n5348);
   U4248 : OAI21_X1 port map( B1 => n6087, B2 => n5868, A => n5349, ZN => n3154
                           );
   U4249 : NAND2_X1 port map( A1 => n1828, A2 => n6871, ZN => n5349);
   U4250 : OAI21_X1 port map( B1 => n6088, B2 => n5869, A => n5350, ZN => n3153
                           );
   U4251 : NAND2_X1 port map( A1 => n1828, A2 => n6868, ZN => n5350);
   U4252 : OAI21_X1 port map( B1 => n6089, B2 => n5868, A => n5351, ZN => n3152
                           );
   U4253 : NAND2_X1 port map( A1 => n1828, A2 => n6865, ZN => n5351);
   U4254 : OAI21_X1 port map( B1 => n6090, B2 => n5868, A => n5352, ZN => n3151
                           );
   U4255 : NAND2_X1 port map( A1 => n1828, A2 => n6862, ZN => n5352);
   U4256 : NAND2_X1 port map( A1 => n1692, A2 => n1590, ZN => n1828);
   U4258 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n6050, ZN => n5353);
   U4259 : NOR2_X1 port map( A1 => n5354, A2 => n6047, ZN => n1692);
   U4260 : OR2_X1 port map( A1 => ADD_WR(3), A2 => n2273, ZN => n5354);
   U4261 : OAI21_X1 port map( B1 => n6059, B2 => n5355, A => n5356, ZN => n3150
                           );
   U4262 : NAND2_X1 port map( A1 => n5565, A2 => n6937, ZN => n5356);
   U4263 : OAI21_X1 port map( B1 => n6060, B2 => n5567, A => n5357, ZN => n3149
                           );
   U4264 : NAND2_X1 port map( A1 => n5565, A2 => n6935, ZN => n5357);
   U4265 : OAI21_X1 port map( B1 => n6061, B2 => n5355, A => n5358, ZN => n3148
                           );
   U4266 : NAND2_X1 port map( A1 => n5565, A2 => n6933, ZN => n5358);
   U4267 : OAI21_X1 port map( B1 => n6062, B2 => n5567, A => n5359, ZN => n3147
                           );
   U4268 : NAND2_X1 port map( A1 => n5565, A2 => n6931, ZN => n5359);
   U4269 : OAI21_X1 port map( B1 => n6063, B2 => n5567, A => n5360, ZN => n3146
                           );
   U4270 : NAND2_X1 port map( A1 => n5565, A2 => n6929, ZN => n5360);
   U4271 : OAI21_X1 port map( B1 => n6064, B2 => n5355, A => n5361, ZN => n3145
                           );
   U4272 : NAND2_X1 port map( A1 => n5567, A2 => n6927, ZN => n5361);
   U4273 : OAI21_X1 port map( B1 => n6065, B2 => n5355, A => n5362, ZN => n3144
                           );
   U4274 : NAND2_X1 port map( A1 => n5565, A2 => n6925, ZN => n5362);
   U4275 : OAI21_X1 port map( B1 => n6066, B2 => n5355, A => n5363, ZN => n3143
                           );
   U4276 : NAND2_X1 port map( A1 => n5567, A2 => n6923, ZN => n5363);
   U4277 : OAI21_X1 port map( B1 => n5481, B2 => n5355, A => n5364, ZN => n3142
                           );
   U4278 : NAND2_X1 port map( A1 => n5567, A2 => n6921, ZN => n5364);
   U4279 : OAI21_X1 port map( B1 => n6068, B2 => n5355, A => n5365, ZN => n3141
                           );
   U4280 : NAND2_X1 port map( A1 => n5567, A2 => n6919, ZN => n5365);
   U4281 : OAI21_X1 port map( B1 => n6069, B2 => n5355, A => n5366, ZN => n3140
                           );
   U4282 : NAND2_X1 port map( A1 => n5567, A2 => n6917, ZN => n5366);
   U4283 : OAI21_X1 port map( B1 => n6070, B2 => n5567, A => n5367, ZN => n3139
                           );
   U4284 : NAND2_X1 port map( A1 => n5567, A2 => n6915, ZN => n5367);
   U4285 : OAI21_X1 port map( B1 => n6071, B2 => n5565, A => n5368, ZN => n3138
                           );
   U4286 : NAND2_X1 port map( A1 => n5567, A2 => n6913, ZN => n5368);
   U4287 : OAI21_X1 port map( B1 => n6072, B2 => n5567, A => n5369, ZN => n3137
                           );
   U4288 : NAND2_X1 port map( A1 => n5565, A2 => n6911, ZN => n5369);
   U4289 : OAI21_X1 port map( B1 => n5499, B2 => n5355, A => n5370, ZN => n3136
                           );
   U4290 : NAND2_X1 port map( A1 => n5567, A2 => n6909, ZN => n5370);
   U4291 : OAI21_X1 port map( B1 => n6074, B2 => n5567, A => n5371, ZN => n3135
                           );
   U4292 : NAND2_X1 port map( A1 => n5567, A2 => n6907, ZN => n5371);
   U4293 : OAI21_X1 port map( B1 => n6075, B2 => n5355, A => n5372, ZN => n3134
                           );
   U4294 : NAND2_X1 port map( A1 => n5567, A2 => n6905, ZN => n5372);
   U4295 : OAI21_X1 port map( B1 => n6076, B2 => n5355, A => n5373, ZN => n3133
                           );
   U4296 : NAND2_X1 port map( A1 => n5565, A2 => n6902, ZN => n5373);
   U4297 : OAI21_X1 port map( B1 => n6077, B2 => n5355, A => n5374, ZN => n3132
                           );
   U4298 : NAND2_X1 port map( A1 => n5567, A2 => n6899, ZN => n5374);
   U4299 : OAI21_X1 port map( B1 => n6078, B2 => n5355, A => n5375, ZN => n3131
                           );
   U4300 : NAND2_X1 port map( A1 => n5565, A2 => n6896, ZN => n5375);
   U4301 : OAI21_X1 port map( B1 => n6079, B2 => n5355, A => n5376, ZN => n3130
                           );
   U4302 : NAND2_X1 port map( A1 => n5567, A2 => n6893, ZN => n5376);
   U4303 : OAI21_X1 port map( B1 => n6080, B2 => n5355, A => n5377, ZN => n3129
                           );
   U4304 : NAND2_X1 port map( A1 => n5565, A2 => n6890, ZN => n5377);
   U4305 : OAI21_X1 port map( B1 => n5523, B2 => n5355, A => n5378, ZN => n3128
                           );
   U4306 : NAND2_X1 port map( A1 => n5567, A2 => n6887, ZN => n5378);
   U4307 : OAI21_X1 port map( B1 => n6082, B2 => n5355, A => n5379, ZN => n3127
                           );
   U4308 : NAND2_X1 port map( A1 => n5565, A2 => n6884, ZN => n5379);
   U4309 : OAI21_X1 port map( B1 => n6083, B2 => n5355, A => n5380, ZN => n3126
                           );
   U4310 : NAND2_X1 port map( A1 => n5565, A2 => n6881, ZN => n5380);
   U4311 : OAI21_X1 port map( B1 => n6084, B2 => n5355, A => n5381, ZN => n3125
                           );
   U4312 : NAND2_X1 port map( A1 => n5565, A2 => n6878, ZN => n5381);
   U4313 : OAI21_X1 port map( B1 => n6085, B2 => n5355, A => n5382, ZN => n3124
                           );
   U4314 : NAND2_X1 port map( A1 => n5565, A2 => n6875, ZN => n5382);
   U4315 : OAI21_X1 port map( B1 => n6086, B2 => n5355, A => n5383, ZN => n3123
                           );
   U4316 : NAND2_X1 port map( A1 => n5565, A2 => n6872, ZN => n5383);
   U4317 : OAI21_X1 port map( B1 => n6087, B2 => n5355, A => n5384, ZN => n3122
                           );
   U4318 : NAND2_X1 port map( A1 => n5565, A2 => n6869, ZN => n5384);
   U4319 : OAI21_X1 port map( B1 => n6088, B2 => n5355, A => n5385, ZN => n3121
                           );
   U4320 : NAND2_X1 port map( A1 => n5565, A2 => n6866, ZN => n5385);
   U4321 : OAI21_X1 port map( B1 => n6089, B2 => n5355, A => n5386, ZN => n3120
                           );
   U4322 : NAND2_X1 port map( A1 => n5565, A2 => n6863, ZN => n5386);
   U4323 : OAI21_X1 port map( B1 => n6090, B2 => n5567, A => n5387, ZN => n3119
                           );
   U4324 : NAND2_X1 port map( A1 => n5565, A2 => n6860, ZN => n5387);
   U4325 : NAND2_X1 port map( A1 => n1777, A2 => n1521, ZN => n5355);
   U4326 : NOR2_X1 port map( A1 => n5388, A2 => n6049, ZN => n1521);
   U4327 : OR2_X1 port map( A1 => ADD_WR(1), A2 => n6050, ZN => n5388);
   U4328 : OAI21_X1 port map( B1 => n6059, B2 => n5562, A => n5390, ZN => n3118
                           );
   U4329 : NAND2_X1 port map( A1 => n5389, A2 => n6938, ZN => n5390);
   U4330 : OAI21_X1 port map( B1 => n6060, B2 => n5564, A => n5391, ZN => n3117
                           );
   U4331 : NAND2_X1 port map( A1 => n5389, A2 => n6936, ZN => n5391);
   U4332 : OAI21_X1 port map( B1 => n6061, B2 => n5562, A => n5392, ZN => n3116
                           );
   U4333 : NAND2_X1 port map( A1 => n5389, A2 => n6934, ZN => n5392);
   U4334 : OAI21_X1 port map( B1 => n6062, B2 => n5562, A => n5393, ZN => n3115
                           );
   U4335 : NAND2_X1 port map( A1 => n5389, A2 => n6932, ZN => n5393);
   U4336 : OAI21_X1 port map( B1 => n6063, B2 => n5564, A => n5394, ZN => n3114
                           );
   U4337 : NAND2_X1 port map( A1 => n5564, A2 => n6930, ZN => n5394);
   U4338 : OAI21_X1 port map( B1 => n6064, B2 => n5562, A => n5395, ZN => n3113
                           );
   U4339 : NAND2_X1 port map( A1 => n5389, A2 => n6928, ZN => n5395);
   U4340 : OAI21_X1 port map( B1 => n6065, B2 => n5562, A => n5396, ZN => n3112
                           );
   U4341 : NAND2_X1 port map( A1 => n5389, A2 => n6926, ZN => n5396);
   U4342 : OAI21_X1 port map( B1 => n6066, B2 => n5562, A => n5397, ZN => n3111
                           );
   U4343 : NAND2_X1 port map( A1 => n5562, A2 => n6924, ZN => n5397);
   U4344 : OAI21_X1 port map( B1 => n5481, B2 => n5562, A => n5398, ZN => n3110
                           );
   U4345 : NAND2_X1 port map( A1 => n5389, A2 => n6922, ZN => n5398);
   U4346 : OAI21_X1 port map( B1 => n6068, B2 => n5562, A => n5399, ZN => n3109
                           );
   U4347 : NAND2_X1 port map( A1 => n5389, A2 => n6920, ZN => n5399);
   U4348 : OAI21_X1 port map( B1 => n6069, B2 => n5562, A => n5400, ZN => n3108
                           );
   U4349 : NAND2_X1 port map( A1 => n5389, A2 => n6918, ZN => n5400);
   U4350 : OAI21_X1 port map( B1 => n6070, B2 => n5562, A => n5401, ZN => n3107
                           );
   U4351 : NAND2_X1 port map( A1 => n5389, A2 => n6916, ZN => n5401);
   U4352 : OAI21_X1 port map( B1 => n6071, B2 => n5562, A => n5402, ZN => n3106
                           );
   U4353 : NAND2_X1 port map( A1 => n5389, A2 => n6914, ZN => n5402);
   U4354 : OAI21_X1 port map( B1 => n6072, B2 => n5562, A => n5403, ZN => n3105
                           );
   U4355 : NAND2_X1 port map( A1 => n5389, A2 => n6912, ZN => n5403);
   U4356 : OAI21_X1 port map( B1 => n5499, B2 => n5562, A => n5404, ZN => n3104
                           );
   U4357 : NAND2_X1 port map( A1 => n5389, A2 => n6910, ZN => n5404);
   U4358 : OAI21_X1 port map( B1 => n6074, B2 => n5564, A => n5405, ZN => n3103
                           );
   U4359 : NAND2_X1 port map( A1 => n5389, A2 => n6908, ZN => n5405);
   U4360 : OAI21_X1 port map( B1 => n6075, B2 => n5562, A => n5406, ZN => n3102
                           );
   U4361 : NAND2_X1 port map( A1 => n5389, A2 => n6906, ZN => n5406);
   U4362 : OAI21_X1 port map( B1 => n6076, B2 => n5564, A => n5407, ZN => n3101
                           );
   U4363 : NAND2_X1 port map( A1 => n5564, A2 => n6903, ZN => n5407);
   U4364 : OAI21_X1 port map( B1 => n6077, B2 => n5562, A => n5408, ZN => n3100
                           );
   U4365 : NAND2_X1 port map( A1 => n5564, A2 => n6900, ZN => n5408);
   U4366 : OAI21_X1 port map( B1 => n6078, B2 => n5564, A => n5409, ZN => n3099
                           );
   U4367 : NAND2_X1 port map( A1 => n5564, A2 => n6897, ZN => n5409);
   U4368 : OAI21_X1 port map( B1 => n6079, B2 => n5562, A => n5410, ZN => n3098
                           );
   U4369 : NAND2_X1 port map( A1 => n5564, A2 => n6894, ZN => n5410);
   U4370 : OAI21_X1 port map( B1 => n6080, B2 => n5564, A => n5411, ZN => n3097
                           );
   U4371 : NAND2_X1 port map( A1 => n5564, A2 => n6891, ZN => n5411);
   U4372 : OAI21_X1 port map( B1 => n5523, B2 => n5562, A => n5412, ZN => n3096
                           );
   U4373 : NAND2_X1 port map( A1 => n5564, A2 => n6888, ZN => n5412);
   U4374 : OAI21_X1 port map( B1 => n6082, B2 => n5564, A => n5413, ZN => n3095
                           );
   U4375 : NAND2_X1 port map( A1 => n5564, A2 => n6885, ZN => n5413);
   U4376 : OAI21_X1 port map( B1 => n6083, B2 => n5562, A => n5414, ZN => n3094
                           );
   U4377 : NAND2_X1 port map( A1 => n5389, A2 => n6882, ZN => n5414);
   U4378 : OAI21_X1 port map( B1 => n6084, B2 => n5389, A => n5415, ZN => n3093
                           );
   U4379 : NAND2_X1 port map( A1 => n5389, A2 => n6879, ZN => n5415);
   U4380 : OAI21_X1 port map( B1 => n6085, B2 => n5564, A => n5416, ZN => n3092
                           );
   U4381 : NAND2_X1 port map( A1 => n5389, A2 => n6876, ZN => n5416);
   U4382 : OAI21_X1 port map( B1 => n6086, B2 => n5564, A => n5417, ZN => n3091
                           );
   U4383 : NAND2_X1 port map( A1 => n5389, A2 => n6873, ZN => n5417);
   U4384 : OAI21_X1 port map( B1 => n6087, B2 => n5564, A => n5418, ZN => n3090
                           );
   U4385 : NAND2_X1 port map( A1 => n5389, A2 => n6870, ZN => n5418);
   U4386 : OAI21_X1 port map( B1 => n6088, B2 => n5564, A => n5419, ZN => n3089
                           );
   U4387 : NAND2_X1 port map( A1 => n5389, A2 => n6867, ZN => n5419);
   U4388 : OAI21_X1 port map( B1 => n6089, B2 => n5564, A => n5420, ZN => n3088
                           );
   U4389 : NAND2_X1 port map( A1 => n5389, A2 => n6864, ZN => n5420);
   U4390 : OAI21_X1 port map( B1 => n6090, B2 => n5562, A => n5421, ZN => n3087
                           );
   U4391 : NAND2_X1 port map( A1 => n5389, A2 => n6861, ZN => n5421);
   U4392 : NAND2_X1 port map( A1 => n2110, A2 => n1777, ZN => n5389);
   U4393 : NOR2_X1 port map( A1 => n5422, A2 => n6047, ZN => n1777);
   U4394 : OR2_X1 port map( A1 => n2273, A2 => n6048, ZN => n5422);
   U4395 : NOR2_X1 port map( A1 => n2453, A2 => ADD_WR(0), ZN => n2110);
   U4396 : OR2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n2453);
   U4397 : OAI21_X1 port map( B1 => n6059, B2 => n5556, A => n5424, ZN => n3086
                           );
   U4398 : NAND2_X1 port map( A1 => n5423, A2 => n6667, ZN => n5424);
   U4399 : OAI21_X1 port map( B1 => n6060, B2 => n5557, A => n5425, ZN => n3085
                           );
   U4400 : NAND2_X1 port map( A1 => n5423, A2 => n6666, ZN => n5425);
   U4401 : OAI21_X1 port map( B1 => n6061, B2 => n5556, A => n5426, ZN => n3084
                           );
   U4402 : NAND2_X1 port map( A1 => n5423, A2 => n6665, ZN => n5426);
   U4403 : OAI21_X1 port map( B1 => n6062, B2 => n5556, A => n5427, ZN => n3083
                           );
   U4404 : NAND2_X1 port map( A1 => n5423, A2 => n6664, ZN => n5427);
   U4405 : OAI21_X1 port map( B1 => n6063, B2 => n5557, A => n5428, ZN => n3082
                           );
   U4406 : NAND2_X1 port map( A1 => n5423, A2 => n6663, ZN => n5428);
   U4407 : OAI21_X1 port map( B1 => n6064, B2 => n5556, A => n5429, ZN => n3081
                           );
   U4408 : NAND2_X1 port map( A1 => n5423, A2 => n6662, ZN => n5429);
   U4409 : OAI21_X1 port map( B1 => n6065, B2 => n5556, A => n5430, ZN => n3080
                           );
   U4410 : NAND2_X1 port map( A1 => n5423, A2 => n6661, ZN => n5430);
   U4411 : OAI21_X1 port map( B1 => n6066, B2 => n5556, A => n5431, ZN => n3079
                           );
   U4412 : NAND2_X1 port map( A1 => n5557, A2 => n6660, ZN => n5431);
   U4413 : OAI21_X1 port map( B1 => n5481, B2 => n5556, A => n5432, ZN => n3078
                           );
   U4414 : NAND2_X1 port map( A1 => n5556, A2 => n6659, ZN => n5432);
   U4415 : OAI21_X1 port map( B1 => n6068, B2 => n5556, A => n5433, ZN => n3077
                           );
   U4416 : NAND2_X1 port map( A1 => n5557, A2 => n6658, ZN => n5433);
   U4417 : OAI21_X1 port map( B1 => n6069, B2 => n5556, A => n5434, ZN => n3076
                           );
   U4418 : NAND2_X1 port map( A1 => n5556, A2 => n6657, ZN => n5434);
   U4419 : OAI21_X1 port map( B1 => n6070, B2 => n5556, A => n5435, ZN => n3075
                           );
   U4420 : NAND2_X1 port map( A1 => n5557, A2 => n6656, ZN => n5435);
   U4421 : OAI21_X1 port map( B1 => n6071, B2 => n5556, A => n5436, ZN => n3074
                           );
   U4422 : NAND2_X1 port map( A1 => n5556, A2 => n6655, ZN => n5436);
   U4423 : OAI21_X1 port map( B1 => n6072, B2 => n5556, A => n5437, ZN => n3073
                           );
   U4424 : NAND2_X1 port map( A1 => n5423, A2 => n6654, ZN => n5437);
   U4425 : OAI21_X1 port map( B1 => n5499, B2 => n5556, A => n5438, ZN => n3072
                           );
   U4426 : NAND2_X1 port map( A1 => n5557, A2 => n6653, ZN => n5438);
   U4427 : OAI21_X1 port map( B1 => n6074, B2 => n5557, A => n5439, ZN => n3071
                           );
   U4428 : NAND2_X1 port map( A1 => n5556, A2 => n6652, ZN => n5439);
   U4429 : OAI21_X1 port map( B1 => n5506, B2 => n5557, A => n5440, ZN => n3070
                           );
   U4430 : NAND2_X1 port map( A1 => n5423, A2 => n6651, ZN => n5440);
   U4431 : OAI21_X1 port map( B1 => n6076, B2 => n5557, A => n5441, ZN => n3069
                           );
   U4432 : NAND2_X1 port map( A1 => n5423, A2 => n6650, ZN => n5441);
   U4433 : OAI21_X1 port map( B1 => n6077, B2 => n5557, A => n5442, ZN => n3068
                           );
   U4434 : NAND2_X1 port map( A1 => n5423, A2 => n6649, ZN => n5442);
   U4435 : OAI21_X1 port map( B1 => n6078, B2 => n5557, A => n5443, ZN => n3067
                           );
   U4436 : NAND2_X1 port map( A1 => n5423, A2 => n6648, ZN => n5443);
   U4437 : OAI21_X1 port map( B1 => n6079, B2 => n5557, A => n5444, ZN => n3066
                           );
   U4438 : NAND2_X1 port map( A1 => n5423, A2 => n6647, ZN => n5444);
   U4439 : OAI21_X1 port map( B1 => n6080, B2 => n5557, A => n5445, ZN => n3065
                           );
   U4440 : NAND2_X1 port map( A1 => n5423, A2 => n6646, ZN => n5445);
   U4441 : OAI21_X1 port map( B1 => n5523, B2 => n5557, A => n5446, ZN => n3064
                           );
   U4442 : NAND2_X1 port map( A1 => n5423, A2 => n6645, ZN => n5446);
   U4443 : OAI21_X1 port map( B1 => n6082, B2 => n5557, A => n5447, ZN => n3063
                           );
   U4444 : NAND2_X1 port map( A1 => n5423, A2 => n6644, ZN => n5447);
   U4445 : OAI21_X1 port map( B1 => n6083, B2 => n5557, A => n5448, ZN => n3062
                           );
   U4446 : NAND2_X1 port map( A1 => n5423, A2 => n6643, ZN => n5448);
   U4447 : OAI21_X1 port map( B1 => n6084, B2 => n5557, A => n5449, ZN => n3061
                           );
   U4448 : NAND2_X1 port map( A1 => n5423, A2 => n6642, ZN => n5449);
   U4449 : OAI21_X1 port map( B1 => n6085, B2 => n5557, A => n5450, ZN => n3060
                           );
   U4450 : NAND2_X1 port map( A1 => n5423, A2 => n6641, ZN => n5450);
   U4451 : OAI21_X1 port map( B1 => n6086, B2 => n5557, A => n5451, ZN => n3059
                           );
   U4452 : NAND2_X1 port map( A1 => n5423, A2 => n6640, ZN => n5451);
   U4453 : OAI21_X1 port map( B1 => n6087, B2 => n5556, A => n5452, ZN => n3058
                           );
   U4454 : NAND2_X1 port map( A1 => n5423, A2 => n6639, ZN => n5452);
   U4455 : OAI21_X1 port map( B1 => n6088, B2 => n5557, A => n5453, ZN => n3057
                           );
   U4456 : NAND2_X1 port map( A1 => n5423, A2 => n6638, ZN => n5453);
   U4457 : OAI21_X1 port map( B1 => n6089, B2 => n5556, A => n5454, ZN => n3056
                           );
   U4458 : NAND2_X1 port map( A1 => n5423, A2 => n6637, ZN => n5454);
   U4459 : OAI21_X1 port map( B1 => n6090, B2 => n5556, A => n5455, ZN => n3055
                           );
   U4460 : NAND2_X1 port map( A1 => n5423, A2 => n6636, ZN => n5455);
   U4461 : NAND2_X1 port map( A1 => n1812, A2 => n1520, ZN => n5423);
   U4462 : NOR3_X1 port map( A1 => n2273, A2 => ADD_WR(4), A3 => ADD_WR(3), ZN 
                           => n1520);
   U4463 : NAND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n2273);
   U4464 : NOR2_X1 port map( A1 => n5456, A2 => n6049, ZN => n1812);
   U4465 : OR2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n5456);
   U20 : CLKBUF_X1 port map( A => n2342, Z => n5775);
   U21 : CLKBUF_X1 port map( A => n2420, Z => n5764);
   U24 : CLKBUF_X1 port map( A => n2011, Z => n5829);
   U25 : CLKBUF_X1 port map( A => n2077, Z => n5818);
   U34 : CLKBUF_X1 port map( A => n2231, Z => n5793);
   U37 : CLKBUF_X1 port map( A => n1879, Z => n5854);
   U47 : CLKBUF_X1 port map( A => n1487, Z => n5925);
   U52 : CLKBUF_X1 port map( A => n2342, Z => n5777);
   U54 : CLKBUF_X1 port map( A => n2011, Z => n5831);
   U58 : CLKBUF_X1 port map( A => n2231, Z => n5795);
   U72 : CLKBUF_X1 port map( A => n1779, Z => n5871);
   U79 : CLKBUF_X1 port map( A => n1591, Z => n5907);
   U83 : CLKBUF_X1 port map( A => n5355, Z => n5565);
   U84 : CLKBUF_X1 port map( A => n1693, Z => n5890);
   U92 : CLKBUF_X1 port map( A => n2111, Z => n5812);
   U99 : CLKBUF_X1 port map( A => n1779, Z => n5873);
   U103 : CLKBUF_X1 port map( A => n1591, Z => n5909);
   U105 : CLKBUF_X1 port map( A => n5355, Z => n5567);
   U112 : CLKBUF_X1 port map( A => n2274, Z => n5790);
   U113 : CLKBUF_X1 port map( A => n2274, Z => n5791);
   U115 : CLKBUF_X1 port map( A => n2308, Z => n5785);
   U116 : CLKBUF_X1 port map( A => n5423, Z => n5557);
   U117 : CLKBUF_X1 port map( A => n5423, Z => n5556);
   U121 : CLKBUF_X1 port map( A => n2386, Z => n5773);
   U127 : CLKBUF_X1 port map( A => n5389, Z => n5562);
   U131 : CLKBUF_X1 port map( A => n2044, Z => n5827);
   U135 : CLKBUF_X1 port map( A => n1625, Z => n5904);
   U138 : CLKBUF_X1 port map( A => n2148, Z => n5808);
   U139 : CLKBUF_X1 port map( A => n2148, Z => n5809);
   U141 : CLKBUF_X1 port map( A => n1557, Z => n5916);
   U142 : CLKBUF_X1 port map( A => n1522, Z => n5923);
   U143 : CLKBUF_X1 port map( A => n1522, Z => n5922);
   U145 : CLKBUF_X1 port map( A => n2189, Z => n5803);
   U149 : CLKBUF_X1 port map( A => n1846, Z => n5863);
   U154 : CLKBUF_X1 port map( A => n1912, Z => n5850);
   U155 : CLKBUF_X1 port map( A => n1912, Z => n5851);
   U157 : CLKBUF_X1 port map( A => n1945, Z => n5845);
   U159 : CLKBUF_X1 port map( A => n1744, Z => n5880);
   U162 : CLKBUF_X1 port map( A => n1726, Z => n5887);
   U163 : CLKBUF_X1 port map( A => n1726, Z => n5886);
   U165 : CLKBUF_X1 port map( A => n1978, Z => n5839);
   U166 : CLKBUF_X1 port map( A => n1828, Z => n5869);
   U167 : CLKBUF_X1 port map( A => n1828, Z => n5868);
   U169 : CLKBUF_X1 port map( A => n1659, Z => n5898);
   U202 : CLKBUF_X1 port map( A => n4451, Z => n5649);
   U208 : CLKBUF_X1 port map( A => n2469, Z => n5745);
   U223 : CLKBUF_X1 port map( A => n4490, Z => n5581);
   U228 : CLKBUF_X1 port map( A => n2508, Z => n5677);
   U232 : CLKBUF_X1 port map( A => n4478, Z => n5605);
   U236 : CLKBUF_X1 port map( A => n2496, Z => n5701);
   U243 : CLKBUF_X1 port map( A => n4479, Z => n5601);
   U244 : CLKBUF_X1 port map( A => n4462, Z => n5629);
   U248 : CLKBUF_X1 port map( A => n2497, Z => n5697);
   U249 : CLKBUF_X1 port map( A => n2480, Z => n5725);
   U273 : CLKBUF_X1 port map( A => n4491, Z => n5577);
   U282 : CLKBUF_X1 port map( A => n2509, Z => n5673);
   U305 : CLKBUF_X1 port map( A => n4461, Z => n5633);
   U306 : CLKBUF_X1 port map( A => n4486, Z => n5588);
   U307 : CLKBUF_X1 port map( A => n4492, Z => n5576);
   U308 : CLKBUF_X1 port map( A => n2477, Z => n5735);
   U309 : CLKBUF_X1 port map( A => n2479, Z => n5729);
   U310 : CLKBUF_X1 port map( A => n2493, Z => n5705);
   U311 : CLKBUF_X1 port map( A => n2504, Z => n5684);
   U312 : CLKBUF_X1 port map( A => n2510, Z => n5672);
   U313 : CLKBUF_X1 port map( A => n4447, Z => n5657);
   U314 : CLKBUF_X1 port map( A => n2465, Z => n5753);
   U315 : CLKBUF_X1 port map( A => n4480, Z => n5600);
   U316 : CLKBUF_X1 port map( A => n2498, Z => n5696);
   U317 : CLKBUF_X1 port map( A => n4453, Z => n5645);
   U319 : CLKBUF_X1 port map( A => n4484, Z => n5594);
   U320 : CLKBUF_X1 port map( A => n2471, Z => n5741);
   U322 : CLKBUF_X1 port map( A => n2502, Z => n5690);
   U323 : CLKBUF_X1 port map( A => n4463, Z => n5627);
   U324 : CLKBUF_X1 port map( A => n4473, Z => n5615);
   U325 : CLKBUF_X1 port map( A => n4475, Z => n5609);
   U327 : CLKBUF_X1 port map( A => n2481, Z => n5723);
   U328 : CLKBUF_X1 port map( A => n2491, Z => n5711);
   U330 : CLKBUF_X1 port map( A => n4459, Z => n5639);
   U331 : CLKBUF_X1 port map( A => n4465, Z => n5621);
   U333 : CLKBUF_X1 port map( A => n2483, Z => n5717);
   U335 : CLKBUF_X1 port map( A => n4444, Z => n5663);
   U336 : CLKBUF_X1 port map( A => n2462, Z => n5759);
   U338 : CLKBUF_X1 port map( A => n4454, Z => n5642);
   U342 : CLKBUF_X1 port map( A => n4464, Z => n5624);
   U343 : CLKBUF_X1 port map( A => n4448, Z => n5654);
   U344 : CLKBUF_X1 port map( A => n4474, Z => n5612);
   U345 : CLKBUF_X1 port map( A => n4485, Z => n5591);
   U346 : CLKBUF_X1 port map( A => n4487, Z => n5585);
   U347 : CLKBUF_X1 port map( A => n2466, Z => n5750);
   U348 : CLKBUF_X1 port map( A => n2472, Z => n5738);
   U349 : CLKBUF_X1 port map( A => n2492, Z => n5708);
   U350 : CLKBUF_X1 port map( A => n2503, Z => n5687);
   U351 : CLKBUF_X1 port map( A => n2505, Z => n5681);
   U352 : CLKBUF_X1 port map( A => n4460, Z => n5636);
   U353 : CLKBUF_X1 port map( A => n4466, Z => n5618);
   U355 : CLKBUF_X1 port map( A => n4493, Z => n5573);
   U356 : CLKBUF_X1 port map( A => n2478, Z => n5732);
   U357 : CLKBUF_X1 port map( A => n2482, Z => n5720);
   U358 : CLKBUF_X1 port map( A => n2484, Z => n5714);
   U360 : CLKBUF_X1 port map( A => n2511, Z => n5669);
   U361 : CLKBUF_X1 port map( A => n4452, Z => n5648);
   U362 : CLKBUF_X1 port map( A => n4481, Z => n5597);
   U363 : CLKBUF_X1 port map( A => n2470, Z => n5744);
   U364 : CLKBUF_X1 port map( A => n2499, Z => n5693);
   U365 : CLKBUF_X1 port map( A => n4445, Z => n5660);
   U366 : CLKBUF_X1 port map( A => n2463, Z => n5756);
   U367 : CLKBUF_X1 port map( A => n4442, Z => n5666);
   U368 : CLKBUF_X1 port map( A => n2460, Z => n5762);
   U371 : CLKBUF_X1 port map( A => n6075, Z => n5506);
   U402 : CLKBUF_X1 port map( A => n6076, Z => n5509);
   U412 : CLKBUF_X1 port map( A => n6081, Z => n5523);
   U420 : CLKBUF_X1 port map( A => n6073, Z => n5499);
   U426 : CLKBUF_X1 port map( A => n6067, Z => n5481);
   U435 : CLKBUF_X1 port map( A => n6090, Z => n5552);
   U436 : CLKBUF_X1 port map( A => n6089, Z => n5549);
   U437 : CLKBUF_X1 port map( A => n6088, Z => n5546);
   U438 : CLKBUF_X1 port map( A => n6087, Z => n5543);
   U439 : CLKBUF_X1 port map( A => n6086, Z => n5540);
   U440 : CLKBUF_X1 port map( A => n6085, Z => n5537);
   U441 : CLKBUF_X1 port map( A => n6084, Z => n5534);
   U442 : CLKBUF_X1 port map( A => n6083, Z => n5531);
   U443 : CLKBUF_X1 port map( A => n6082, Z => n5528);
   U445 : CLKBUF_X1 port map( A => n6080, Z => n5522);
   U446 : CLKBUF_X1 port map( A => n6079, Z => n5519);
   U447 : CLKBUF_X1 port map( A => n6078, Z => n5516);
   U448 : CLKBUF_X1 port map( A => n6077, Z => n5513);
   U451 : CLKBUF_X1 port map( A => n6074, Z => n5504);
   U453 : CLKBUF_X1 port map( A => n6072, Z => n5498);
   U454 : CLKBUF_X1 port map( A => n6071, Z => n5495);
   U455 : CLKBUF_X1 port map( A => n6070, Z => n5492);
   U456 : CLKBUF_X1 port map( A => n6069, Z => n5489);
   U457 : CLKBUF_X1 port map( A => n6068, Z => n5486);
   U459 : CLKBUF_X1 port map( A => n6066, Z => n5480);
   U460 : CLKBUF_X1 port map( A => n6065, Z => n5477);
   U461 : CLKBUF_X1 port map( A => n6064, Z => n5474);
   U462 : CLKBUF_X1 port map( A => n6063, Z => n5471);
   U463 : CLKBUF_X1 port map( A => n6062, Z => n5468);
   U464 : CLKBUF_X1 port map( A => n6061, Z => n5465);
   U465 : CLKBUF_X1 port map( A => n6060, Z => n5462);
   U466 : CLKBUF_X1 port map( A => n6059, Z => n5459);
   U467 : INV_X1 port map( A => ADD_WR(2), ZN => n6049);
   U468 : INV_X1 port map( A => ADD_WR(0), ZN => n6050);
   U469 : INV_X1 port map( A => ADD_WR(4), ZN => n6047);
   U470 : INV_X1 port map( A => ADD_WR(3), ZN => n6048);
   U495 : INV_X1 port map( A => ADD_RD2(0), ZN => n6058);
   U496 : INV_X1 port map( A => ADD_RD1(0), ZN => n6054);
   U497 : INV_X1 port map( A => WR, ZN => n6603);
   U506 : INV_X1 port map( A => ADD_RD2(4), ZN => n6055);
   U507 : INV_X1 port map( A => ADD_RD1(4), ZN => n6051);
   U4894 : INV_X1 port map( A => DATAIN(0), ZN => n6090);
   U4895 : INV_X1 port map( A => DATAIN(1), ZN => n6089);
   U4896 : INV_X1 port map( A => DATAIN(2), ZN => n6088);
   U4897 : INV_X1 port map( A => DATAIN(3), ZN => n6087);
   U4898 : INV_X1 port map( A => DATAIN(4), ZN => n6086);
   U4899 : INV_X1 port map( A => DATAIN(5), ZN => n6085);
   U4900 : INV_X1 port map( A => DATAIN(6), ZN => n6084);
   U4901 : INV_X1 port map( A => DATAIN(7), ZN => n6083);
   U4902 : INV_X1 port map( A => DATAIN(8), ZN => n6082);
   U4903 : INV_X1 port map( A => DATAIN(9), ZN => n6081);
   U4904 : INV_X1 port map( A => DATAIN(10), ZN => n6080);
   U4905 : INV_X1 port map( A => DATAIN(11), ZN => n6079);
   U4906 : INV_X1 port map( A => DATAIN(12), ZN => n6078);
   U4907 : INV_X1 port map( A => DATAIN(13), ZN => n6077);
   U4908 : INV_X1 port map( A => DATAIN(14), ZN => n6076);
   U4909 : INV_X1 port map( A => DATAIN(15), ZN => n6075);
   U4910 : INV_X1 port map( A => DATAIN(16), ZN => n6074);
   U4911 : INV_X1 port map( A => DATAIN(17), ZN => n6073);
   U4912 : INV_X1 port map( A => DATAIN(18), ZN => n6072);
   U4913 : INV_X1 port map( A => DATAIN(19), ZN => n6071);
   U4914 : INV_X1 port map( A => DATAIN(20), ZN => n6070);
   U4915 : INV_X1 port map( A => DATAIN(21), ZN => n6069);
   U4916 : INV_X1 port map( A => DATAIN(22), ZN => n6068);
   U4917 : INV_X1 port map( A => DATAIN(23), ZN => n6067);
   U4918 : INV_X1 port map( A => DATAIN(24), ZN => n6066);
   U4919 : INV_X1 port map( A => DATAIN(25), ZN => n6065);
   U4920 : INV_X1 port map( A => DATAIN(26), ZN => n6064);
   U4921 : INV_X1 port map( A => DATAIN(27), ZN => n6063);
   U4922 : INV_X1 port map( A => DATAIN(28), ZN => n6062);
   U4923 : INV_X1 port map( A => DATAIN(29), ZN => n6061);
   U4924 : INV_X1 port map( A => DATAIN(30), ZN => n6060);
   U4925 : INV_X1 port map( A => DATAIN(31), ZN => n6059);
   U4926 : INV_X1 port map( A => ADD_RD2(2), ZN => n6056);
   U4927 : INV_X1 port map( A => ADD_RD2(1), ZN => n6057);
   U4928 : INV_X1 port map( A => ADD_RD1(2), ZN => n6052);
   U4929 : INV_X1 port map( A => ADD_RD1(1), ZN => n6053);
   U4931 : CLKBUF_X1 port map( A => n5389, Z => n5564);
   U4933 : CLKBUF_X1 port map( A => n2420, Z => n5768);
   U4934 : CLKBUF_X1 port map( A => n2386, Z => n5774);
   U4936 : CLKBUF_X1 port map( A => n2308, Z => n5786);
   U4939 : CLKBUF_X1 port map( A => n2189, Z => n5804);
   U4941 : CLKBUF_X1 port map( A => n2111, Z => n5816);
   U4942 : CLKBUF_X1 port map( A => n2077, Z => n5822);
   U4943 : CLKBUF_X1 port map( A => n2044, Z => n5828);
   U4945 : CLKBUF_X1 port map( A => n1978, Z => n5840);
   U4946 : CLKBUF_X1 port map( A => n1945, Z => n5846);
   U4948 : CLKBUF_X1 port map( A => n1879, Z => n5858);
   U4949 : CLKBUF_X1 port map( A => n1846, Z => n5864);
   U4952 : CLKBUF_X1 port map( A => n1744, Z => n5882);
   U4954 : CLKBUF_X1 port map( A => n1693, Z => n5894);
   U4955 : CLKBUF_X1 port map( A => n1659, Z => n5900);
   U4956 : CLKBUF_X1 port map( A => n1625, Z => n5906);
   U4958 : CLKBUF_X1 port map( A => n1557, Z => n5918);
   U4960 : CLKBUF_X1 port map( A => n1487, Z => n5930);
   U4962 : INV_X1 port map( A => ENABLE, ZN => n5932);
   U4964 : INV_X1 port map( A => ENABLE, ZN => n5934);
   U4965 : INV_X1 port map( A => ENABLE, ZN => n5935);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           RESET, Q => n640, QN => n_1073);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           RESET, Q => n639, QN => n_1074);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           RESET, Q => n638, QN => n_1075);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           RESET, Q => n637, QN => n_1076);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           RESET, Q => n636, QN => n_1077);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           RESET, Q => n635, QN => n_1078);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           RESET, Q => n634, QN => n_1079);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           RESET, Q => n633, QN => n_1080);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           RESET, Q => n632, QN => n_1081);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           RESET, Q => n631, QN => n_1082);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           RESET, Q => n630, QN => n_1083);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           RESET, Q => n629, QN => n_1084);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           RESET, Q => n628, QN => n_1085);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           RESET, Q => n627, QN => n_1086);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           RESET, Q => n626, QN => n_1087);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           RESET, Q => n625, QN => n_1088);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           RESET, Q => n624, QN => n_1089);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           RESET, Q => n623, QN => n_1090);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           RESET, Q => n622, QN => n_1091);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           RESET, Q => n621, QN => n_1092);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           RESET, Q => n620, QN => n_1093);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           RESET, Q => n619, QN => n_1094);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           RESET, Q => n618, QN => n_1095);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           RESET, Q => n617, QN => n_1096);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           RESET, Q => n616, QN => n_1097);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           RESET, Q => n615, QN => n_1098);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           RESET, Q => n614, QN => n_1099);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           RESET, Q => n613, QN => n_1100);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           RESET, Q => n612, QN => n_1101);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           RESET, Q => n611, QN => n_1102);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           RESET, Q => n610, QN => n_1103);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           RESET, Q => n609, QN => n_1104);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           RESET, Q => n6939, QN => n_1105);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           RESET, Q => n6940, QN => n_1106);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           RESET, Q => n6941, QN => n_1107);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           RESET, Q => n6942, QN => n_1108);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           RESET, Q => n6943, QN => n_1109);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           RESET, Q => n6944, QN => n_1110);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           RESET, Q => n6945, QN => n_1111);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           RESET, Q => n6946, QN => n_1112);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           RESET, Q => n6947, QN => n_1113);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           RESET, Q => n6948, QN => n_1114);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           RESET, Q => n6949, QN => n_1115);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           RESET, Q => n6950, QN => n_1116);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           RESET, Q => n6951, QN => n_1117);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           RESET, Q => n6952, QN => n_1118);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           RESET, Q => n6953, QN => n_1119);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           RESET, Q => n6954, QN => n_1120);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           RESET, Q => n6955, QN => n_1121);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           RESET, Q => n6956, QN => n_1122);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           RESET, Q => n6957, QN => n_1123);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           RESET, Q => n6958, QN => n_1124);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           RESET, Q => n6959, QN => n_1125);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           RESET, Q => n6960, QN => n_1126);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           RESET, Q => n6961, QN => n_1127);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           RESET, Q => n6962, QN => n_1128);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           RESET, Q => n6963, QN => n_1129);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           RESET, Q => n6964, QN => n_1130);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           RESET, Q => n6965, QN => n_1131);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           RESET, Q => n6966, QN => n_1132);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           RESET, Q => n6967, QN => n_1133);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           RESET, Q => n6968, QN => n_1134);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           RESET, Q => n6969, QN => n_1135);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           RESET, Q => n6970, QN => n_1136);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           RESET, Q => n608, QN => n_1137);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           RESET, Q => n607, QN => n_1138);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           RESET, Q => n606, QN => n_1139);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           RESET, Q => n605, QN => n_1140);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           RESET, Q => n604, QN => n_1141);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           RESET, Q => n603, QN => n_1142);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           RESET, Q => n602, QN => n_1143);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           RESET, Q => n601, QN => n_1144);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           RESET, Q => n600, QN => n_1145);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           RESET, Q => n599, QN => n_1146);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           RESET, Q => n598, QN => n_1147);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           RESET, Q => n597, QN => n_1148);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           RESET, Q => n596, QN => n_1149);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           RESET, Q => n595, QN => n_1150);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           RESET, Q => n594, QN => n_1151);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           RESET, Q => n593, QN => n_1152);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           RESET, Q => n592, QN => n_1153);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           RESET, Q => n591, QN => n_1154);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => 
                           RESET, Q => n590, QN => n_1155);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           RESET, Q => n589, QN => n_1156);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           RESET, Q => n588, QN => n_1157);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           RESET, Q => n587, QN => n_1158);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           RESET, Q => n586, QN => n_1159);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           RESET, Q => n585, QN => n_1160);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           RESET, Q => n584, QN => n_1161);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           RESET, Q => n583, QN => n_1162);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           RESET, Q => n582, QN => n_1163);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           RESET, Q => n581, QN => n_1164);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           RESET, Q => n580, QN => n_1165);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           RESET, Q => n579, QN => n_1166);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           RESET, Q => n578, QN => n_1167);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           RESET, Q => n577, QN => n_1168);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           RESET, Q => n6667, QN => n_1169);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           RESET, Q => n6666, QN => n_1170);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           RESET, Q => n6665, QN => n_1171);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           RESET, Q => n6664, QN => n_1172);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           RESET, Q => n6663, QN => n_1173);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           RESET, Q => n6662, QN => n_1174);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           RESET, Q => n6661, QN => n_1175);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           RESET, Q => n6660, QN => n_1176);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           RESET, Q => n6659, QN => n_1177);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           RESET, Q => n6658, QN => n_1178);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           RESET, Q => n6657, QN => n_1179);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           RESET, Q => n6656, QN => n_1180);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           RESET, Q => n6655, QN => n_1181);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           RESET, Q => n6654, QN => n_1182);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           RESET, Q => n6653, QN => n_1183);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           RESET, Q => n6652, QN => n_1184);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           RESET, Q => n6651, QN => n_1185);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           RESET, Q => n6650, QN => n_1186);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           RESET, Q => n6649, QN => n_1187);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           RESET, Q => n6648, QN => n_1188);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           RESET, Q => n6647, QN => n_1189);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           RESET, Q => n6646, QN => n_1190);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           RESET, Q => n6645, QN => n_1191);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           RESET, Q => n6644, QN => n_1192);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           RESET, Q => n6643, QN => n_1193);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           RESET, Q => n6642, QN => n_1194);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           RESET, Q => n6641, QN => n_1195);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           RESET, Q => n6640, QN => n_1196);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           RESET, Q => n6639, QN => n_1197);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           RESET, Q => n6638, QN => n_1198);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           RESET, Q => n6637, QN => n_1199);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           RESET, Q => n6636, QN => n_1200);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n4189, CK => CLK, RN => 
                           RESET, Q => n7083, QN => n_1201);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n4188, CK => CLK, RN => 
                           RESET, Q => n7082, QN => n_1202);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n4187, CK => CLK, RN => 
                           RESET, Q => n7081, QN => n_1203);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n4186, CK => CLK, RN => 
                           RESET, Q => n7080, QN => n_1204);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n4185, CK => CLK, RN => 
                           RESET, Q => n7079, QN => n_1205);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n4184, CK => CLK, RN => 
                           RESET, Q => n7078, QN => n_1206);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n4183, CK => CLK, RN => 
                           RESET, Q => n7077, QN => n_1207);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n4182, CK => CLK, RN => 
                           RESET, Q => n7076, QN => n_1208);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n4181, CK => CLK, RN => 
                           RESET, Q => n7075, QN => n_1209);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n4180, CK => CLK, RN => 
                           RESET, Q => n7074, QN => n_1210);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n4179, CK => CLK, RN => 
                           RESET, Q => n7073, QN => n_1211);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n4178, CK => CLK, RN => 
                           RESET, Q => n7072, QN => n_1212);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n4177, CK => CLK, RN => 
                           RESET, Q => n7071, QN => n_1213);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n4176, CK => CLK, RN => 
                           RESET, Q => n7070, QN => n_1214);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n4175, CK => CLK, RN => 
                           RESET, Q => n7069, QN => n_1215);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n4174, CK => CLK, RN => 
                           RESET, Q => n7068, QN => n_1216);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n4173, CK => CLK, RN => 
                           RESET, Q => n7067, QN => n_1217);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n4172, CK => CLK, RN => 
                           RESET, Q => n7066, QN => n_1218);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n4171, CK => CLK, RN => 
                           RESET, Q => n7065, QN => n_1219);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n4170, CK => CLK, RN => 
                           RESET, Q => n7064, QN => n_1220);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n4169, CK => CLK, RN => 
                           RESET, Q => n7063, QN => n_1221);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n4168, CK => CLK, RN => 
                           RESET, Q => n7062, QN => n_1222);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n4167, CK => CLK, RN => 
                           RESET, Q => n7061, QN => n_1223);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n4166, CK => CLK, RN => 
                           RESET, Q => n7060, QN => n_1224);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n4165, CK => CLK, RN => 
                           RESET, Q => n7059, QN => n_1225);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n4164, CK => CLK, RN => 
                           RESET, Q => n7058, QN => n_1226);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n4163, CK => CLK, RN => 
                           RESET, Q => n7057, QN => n_1227);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n4162, CK => CLK, RN => 
                           RESET, Q => n7056, QN => n_1228);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n4161, CK => CLK, RN => 
                           RESET, Q => n7055, QN => n_1229);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n4160, CK => CLK, RN => 
                           RESET, Q => n7054, QN => n_1230);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n4159, CK => CLK, RN => 
                           RESET, Q => n7053, QN => n_1231);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n4158, CK => CLK, RN => 
                           RESET, Q => n7052, QN => n_1232);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           RESET, Q => n6764, QN => n_1233);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           RESET, Q => n6765, QN => n_1234);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           RESET, Q => n6766, QN => n_1235);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           RESET, Q => n6767, QN => n_1236);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           RESET, Q => n6768, QN => n_1237);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           RESET, Q => n6769, QN => n_1238);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           RESET, Q => n6770, QN => n_1239);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           RESET, Q => n6771, QN => n_1240);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           RESET, Q => n6772, QN => n_1241);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           RESET, Q => n6773, QN => n_1242);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           RESET, Q => n6774, QN => n_1243);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           RESET, Q => n6775, QN => n_1244);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           RESET, Q => n6776, QN => n_1245);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           RESET, Q => n6777, QN => n_1246);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           RESET, Q => n6778, QN => n_1247);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           RESET, Q => n6779, QN => n_1248);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           RESET, Q => n6780, QN => n_1249);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           RESET, Q => n6781, QN => n_1250);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           RESET, Q => n6782, QN => n_1251);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           RESET, Q => n6783, QN => n_1252);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           RESET, Q => n6784, QN => n_1253);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           RESET, Q => n6785, QN => n_1254);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           RESET, Q => n6786, QN => n_1255);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           RESET, Q => n6787, QN => n_1256);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           RESET, Q => n6788, QN => n_1257);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           RESET, Q => n6789, QN => n_1258);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           RESET, Q => n6790, QN => n_1259);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           RESET, Q => n6791, QN => n_1260);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           RESET, Q => n6792, QN => n_1261);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           RESET, Q => n6793, QN => n_1262);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           RESET, Q => n6794, QN => n_1263);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           RESET, Q => n6795, QN => n_1264);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           RESET, Q => n480, QN => n_1265);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           RESET, Q => n479, QN => n_1266);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           RESET, Q => n478, QN => n_1267);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           RESET, Q => n477, QN => n_1268);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           RESET, Q => n476, QN => n_1269);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           RESET, Q => n475, QN => n_1270);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           RESET, Q => n474, QN => n_1271);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           RESET, Q => n473, QN => n_1272);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           RESET, Q => n472, QN => n_1273);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           RESET, Q => n471, QN => n_1274);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           RESET, Q => n470, QN => n_1275);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           RESET, Q => n469, QN => n_1276);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           RESET, Q => n468, QN => n_1277);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           RESET, Q => n467, QN => n_1278);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           RESET, Q => n466, QN => n_1279);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           RESET, Q => n465, QN => n_1280);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           RESET, Q => n464, QN => n_1281);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           RESET, Q => n463, QN => n_1282);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           RESET, Q => n462, QN => n_1283);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           RESET, Q => n461, QN => n_1284);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           RESET, Q => n460, QN => n_1285);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           RESET, Q => n459, QN => n_1286);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           RESET, Q => n458, QN => n_1287);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           RESET, Q => n457, QN => n_1288);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           RESET, Q => n456, QN => n_1289);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           RESET, Q => n455, QN => n_1290);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           RESET, Q => n454, QN => n_1291);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           RESET, Q => n453, QN => n_1292);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           RESET, Q => n452, QN => n_1293);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           RESET, Q => n451, QN => n_1294);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           RESET, Q => n450, QN => n_1295);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           RESET, Q => n449, QN => n_1296);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           RESET, Q => n576, QN => n_1297);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           RESET, Q => n575, QN => n_1298);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           RESET, Q => n574, QN => n_1299);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           RESET, Q => n573, QN => n_1300);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           RESET, Q => n572, QN => n_1301);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           RESET, Q => n571, QN => n_1302);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           RESET, Q => n570, QN => n_1303);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           RESET, Q => n569, QN => n_1304);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           RESET, Q => n568, QN => n_1305);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           RESET, Q => n567, QN => n_1306);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           RESET, Q => n566, QN => n_1307);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           RESET, Q => n565, QN => n_1308);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           RESET, Q => n564, QN => n_1309);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           RESET, Q => n563, QN => n_1310);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           RESET, Q => n562, QN => n_1311);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           RESET, Q => n561, QN => n_1312);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           RESET, Q => n560, QN => n_1313);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           RESET, Q => n559, QN => n_1314);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           RESET, Q => n558, QN => n_1315);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           RESET, Q => n557, QN => n_1316);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           RESET, Q => n556, QN => n_1317);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           RESET, Q => n555, QN => n_1318);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           RESET, Q => n554, QN => n_1319);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           RESET, Q => n553, QN => n_1320);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           RESET, Q => n552, QN => n_1321);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           RESET, Q => n551, QN => n_1322);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           RESET, Q => n550, QN => n_1323);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           RESET, Q => n549, QN => n_1324);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           RESET, Q => n548, QN => n_1325);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           RESET, Q => n547, QN => n_1326);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           RESET, Q => n546, QN => n_1327);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           RESET, Q => n545, QN => n_1328);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n3422, CK => CLK, RN => 
                           RESET, Q => n448, QN => n_1329);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n3423, CK => CLK, RN => 
                           RESET, Q => n447, QN => n_1330);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n3424, CK => CLK, RN => 
                           RESET, Q => n446, QN => n_1331);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n3425, CK => CLK, RN => 
                           RESET, Q => n445, QN => n_1332);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n3426, CK => CLK, RN => 
                           RESET, Q => n444, QN => n_1333);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n3427, CK => CLK, RN => 
                           RESET, Q => n443, QN => n_1334);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n3428, CK => CLK, RN => 
                           RESET, Q => n442, QN => n_1335);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n3429, CK => CLK, RN => 
                           RESET, Q => n441, QN => n_1336);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n3430, CK => CLK, RN => 
                           RESET, Q => n440, QN => n_1337);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n3431, CK => CLK, RN => 
                           RESET, Q => n439, QN => n_1338);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n3432, CK => CLK, RN => 
                           RESET, Q => n438, QN => n_1339);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n3433, CK => CLK, RN => 
                           RESET, Q => n437, QN => n_1340);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n3434, CK => CLK, RN => 
                           RESET, Q => n436, QN => n_1341);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n3435, CK => CLK, RN => 
                           RESET, Q => n435, QN => n_1342);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n3436, CK => CLK, RN => 
                           RESET, Q => n434, QN => n_1343);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n3437, CK => CLK, RN => 
                           RESET, Q => n433, QN => n_1344);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n3438, CK => CLK, RN => 
                           RESET, Q => n432, QN => n_1345);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n3439, CK => CLK, RN => 
                           RESET, Q => n431, QN => n_1346);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n3440, CK => CLK, RN => 
                           RESET, Q => n430, QN => n_1347);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n3441, CK => CLK, RN => 
                           RESET, Q => n429, QN => n_1348);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n3442, CK => CLK, RN => 
                           RESET, Q => n428, QN => n_1349);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n3443, CK => CLK, RN => 
                           RESET, Q => n427, QN => n_1350);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n3444, CK => CLK, RN => 
                           RESET, Q => n426, QN => n_1351);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n3445, CK => CLK, RN => 
                           RESET, Q => n425, QN => n_1352);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n3446, CK => CLK, RN => 
                           RESET, Q => n424, QN => n_1353);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n3447, CK => CLK, RN => 
                           RESET, Q => n423, QN => n_1354);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n3448, CK => CLK, RN => 
                           RESET, Q => n422, QN => n_1355);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n3449, CK => CLK, RN => 
                           RESET, Q => n421, QN => n_1356);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n3450, CK => CLK, RN => 
                           RESET, Q => n420, QN => n_1357);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n3451, CK => CLK, RN => 
                           RESET, Q => n419, QN => n_1358);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n3452, CK => CLK, RN => 
                           RESET, Q => n418, QN => n_1359);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n3453, CK => CLK, RN => 
                           RESET, Q => n417, QN => n_1360);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n4157, CK => CLK, RN => 
                           RESET, Q => n6710, QN => n_1361);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n4156, CK => CLK, RN => 
                           RESET, Q => n6709, QN => n_1362);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n4155, CK => CLK, RN => 
                           RESET, Q => n6708, QN => n_1363);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n4154, CK => CLK, RN => 
                           RESET, Q => n2270, QN => n_1364);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n4153, CK => CLK, RN => 
                           RESET, Q => n2265, QN => n_1365);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n4152, CK => CLK, RN => 
                           RESET, Q => n2260, QN => n_1366);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n4151, CK => CLK, RN => 
                           RESET, Q => n2255, QN => n_1367);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n4150, CK => CLK, RN => 
                           RESET, Q => n2250, QN => n_1368);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n4149, CK => CLK, RN => 
                           RESET, Q => n2245, QN => n_1369);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n4148, CK => CLK, RN => 
                           RESET, Q => n2240, QN => n_1370);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n4147, CK => CLK, RN => 
                           RESET, Q => n2235, QN => n_1371);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n4146, CK => CLK, RN => 
                           RESET, Q => n2230, QN => n_1372);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n4145, CK => CLK, RN => 
                           RESET, Q => n2225, QN => n_1373);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n4144, CK => CLK, RN => 
                           RESET, Q => n2220, QN => n_1374);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n4143, CK => CLK, RN => 
                           RESET, Q => n2215, QN => n_1375);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n4142, CK => CLK, RN => 
                           RESET, Q => n2210, QN => n_1376);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n4141, CK => CLK, RN => 
                           RESET, Q => n2205, QN => n_1377);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n4140, CK => CLK, RN => 
                           RESET, Q => n2200, QN => n_1378);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n4139, CK => CLK, RN => 
                           RESET, Q => n2195, QN => n_1379);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n4138, CK => CLK, RN => 
                           RESET, Q => n2190, QN => n_1380);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n4137, CK => CLK, RN => 
                           RESET, Q => n2185, QN => n_1381);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n4136, CK => CLK, RN => 
                           RESET, Q => n2180, QN => n_1382);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n4135, CK => CLK, RN => 
                           RESET, Q => n2175, QN => n_1383);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n4134, CK => CLK, RN => 
                           RESET, Q => n2170, QN => n_1384);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n4133, CK => CLK, RN => 
                           RESET, Q => n2165, QN => n_1385);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n4132, CK => CLK, RN => 
                           RESET, Q => n2160, QN => n_1386);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n4131, CK => CLK, RN => 
                           RESET, Q => n2155, QN => n_1387);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n4130, CK => CLK, RN => 
                           RESET, Q => n2150, QN => n_1388);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n4129, CK => CLK, RN => 
                           RESET, Q => n2145, QN => n_1389);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n4128, CK => CLK, RN => 
                           RESET, Q => n2140, QN => n_1390);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n4127, CK => CLK, RN => 
                           RESET, Q => n2135, QN => n_1391);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n4126, CK => CLK, RN => 
                           RESET, Q => n2130, QN => n_1392);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n4125, CK => CLK, RN => 
                           RESET, Q => n7051, QN => n_1393);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n4124, CK => CLK, RN => 
                           RESET, Q => n7050, QN => n_1394);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n4123, CK => CLK, RN => 
                           RESET, Q => n7049, QN => n_1395);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n4122, CK => CLK, RN => 
                           RESET, Q => n7048, QN => n_1396);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n4121, CK => CLK, RN => 
                           RESET, Q => n7047, QN => n_1397);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n4120, CK => CLK, RN => 
                           RESET, Q => n7046, QN => n_1398);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n4119, CK => CLK, RN => 
                           RESET, Q => n7045, QN => n_1399);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n4118, CK => CLK, RN => 
                           RESET, Q => n7044, QN => n_1400);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n4117, CK => CLK, RN => 
                           RESET, Q => n7043, QN => n_1401);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n4116, CK => CLK, RN => 
                           RESET, Q => n7042, QN => n_1402);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n4115, CK => CLK, RN => 
                           RESET, Q => n7041, QN => n_1403);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n4114, CK => CLK, RN => 
                           RESET, Q => n7040, QN => n_1404);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n4113, CK => CLK, RN => 
                           RESET, Q => n7039, QN => n_1405);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n4112, CK => CLK, RN => 
                           RESET, Q => n7038, QN => n_1406);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n4111, CK => CLK, RN => 
                           RESET, Q => n7037, QN => n_1407);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n4110, CK => CLK, RN => 
                           RESET, Q => n7036, QN => n_1408);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n4109, CK => CLK, RN => 
                           RESET, Q => n7035, QN => n_1409);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n4108, CK => CLK, RN => 
                           RESET, Q => n7034, QN => n_1410);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n4107, CK => CLK, RN => 
                           RESET, Q => n7033, QN => n_1411);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n4106, CK => CLK, RN => 
                           RESET, Q => n7032, QN => n_1412);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n4105, CK => CLK, RN => 
                           RESET, Q => n7031, QN => n_1413);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n4104, CK => CLK, RN => 
                           RESET, Q => n7030, QN => n_1414);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n4103, CK => CLK, RN => 
                           RESET, Q => n7029, QN => n_1415);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n4102, CK => CLK, RN => 
                           RESET, Q => n7028, QN => n_1416);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n4101, CK => CLK, RN => 
                           RESET, Q => n7027, QN => n_1417);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n4100, CK => CLK, RN => 
                           RESET, Q => n7026, QN => n_1418);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n4099, CK => CLK, RN => 
                           RESET, Q => n7025, QN => n_1419);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n4098, CK => CLK, RN => 
                           RESET, Q => n7024, QN => n_1420);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n4097, CK => CLK, RN => 
                           RESET, Q => n7023, QN => n_1421);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n4096, CK => CLK, RN => 
                           RESET, Q => n7022, QN => n_1422);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n4095, CK => CLK, RN => 
                           RESET, Q => n7021, QN => n_1423);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n4094, CK => CLK, RN => 
                           RESET, Q => n7020, QN => n_1424);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n3454, CK => CLK, RN => 
                           RESET, Q => n416, QN => n_1425);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n3455, CK => CLK, RN => 
                           RESET, Q => n415, QN => n_1426);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n3456, CK => CLK, RN => 
                           RESET, Q => n414, QN => n_1427);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n3457, CK => CLK, RN => 
                           RESET, Q => n413, QN => n_1428);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n3458, CK => CLK, RN => 
                           RESET, Q => n412, QN => n_1429);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n3459, CK => CLK, RN => 
                           RESET, Q => n411, QN => n_1430);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n3460, CK => CLK, RN => 
                           RESET, Q => n410, QN => n_1431);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n3461, CK => CLK, RN => 
                           RESET, Q => n409, QN => n_1432);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n3462, CK => CLK, RN => 
                           RESET, Q => n408, QN => n_1433);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n3463, CK => CLK, RN => 
                           RESET, Q => n407, QN => n_1434);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n3464, CK => CLK, RN => 
                           RESET, Q => n406, QN => n_1435);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n3465, CK => CLK, RN => 
                           RESET, Q => n405, QN => n_1436);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n3466, CK => CLK, RN => 
                           RESET, Q => n404, QN => n_1437);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n3467, CK => CLK, RN => 
                           RESET, Q => n403, QN => n_1438);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n3468, CK => CLK, RN => 
                           RESET, Q => n402, QN => n_1439);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n3469, CK => CLK, RN => 
                           RESET, Q => n401, QN => n_1440);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n3470, CK => CLK, RN => 
                           RESET, Q => n400, QN => n_1441);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n3471, CK => CLK, RN => 
                           RESET, Q => n399, QN => n_1442);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n3472, CK => CLK, RN => 
                           RESET, Q => n398, QN => n_1443);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n3473, CK => CLK, RN => 
                           RESET, Q => n397, QN => n_1444);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n3474, CK => CLK, RN => 
                           RESET, Q => n396, QN => n_1445);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n3475, CK => CLK, RN => 
                           RESET, Q => n395, QN => n_1446);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n3476, CK => CLK, RN => 
                           RESET, Q => n394, QN => n_1447);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n3477, CK => CLK, RN => 
                           RESET, Q => n393, QN => n_1448);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n3478, CK => CLK, RN => 
                           RESET, Q => n392, QN => n_1449);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n3479, CK => CLK, RN => 
                           RESET, Q => n391, QN => n_1450);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n3480, CK => CLK, RN => 
                           RESET, Q => n390, QN => n_1451);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n3481, CK => CLK, RN => 
                           RESET, Q => n389, QN => n_1452);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n3482, CK => CLK, RN => 
                           RESET, Q => n388, QN => n_1453);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n3483, CK => CLK, RN => 
                           RESET, Q => n387, QN => n_1454);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n3484, CK => CLK, RN => 
                           RESET, Q => n386, QN => n_1455);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n3485, CK => CLK, RN => 
                           RESET, Q => n385, QN => n_1456);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n3486, CK => CLK, RN => 
                           RESET, Q => n6796, QN => n_1457);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n3487, CK => CLK, RN => 
                           RESET, Q => n6797, QN => n_1458);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n3488, CK => CLK, RN => 
                           RESET, Q => n6798, QN => n_1459);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n3489, CK => CLK, RN => 
                           RESET, Q => n6799, QN => n_1460);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n3490, CK => CLK, RN => 
                           RESET, Q => n6800, QN => n_1461);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n3491, CK => CLK, RN => 
                           RESET, Q => n6801, QN => n_1462);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n3492, CK => CLK, RN => 
                           RESET, Q => n6802, QN => n_1463);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n3493, CK => CLK, RN => 
                           RESET, Q => n6803, QN => n_1464);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n3494, CK => CLK, RN => 
                           RESET, Q => n6804, QN => n_1465);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n3495, CK => CLK, RN => 
                           RESET, Q => n6805, QN => n_1466);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n3496, CK => CLK, RN => 
                           RESET, Q => n6806, QN => n_1467);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n3497, CK => CLK, RN => 
                           RESET, Q => n6807, QN => n_1468);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n3498, CK => CLK, RN => 
                           RESET, Q => n6808, QN => n_1469);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n3499, CK => CLK, RN => 
                           RESET, Q => n6809, QN => n_1470);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n3500, CK => CLK, RN => 
                           RESET, Q => n6810, QN => n_1471);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n3501, CK => CLK, RN => 
                           RESET, Q => n6811, QN => n_1472);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n3502, CK => CLK, RN => 
                           RESET, Q => n6812, QN => n_1473);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n3503, CK => CLK, RN => 
                           RESET, Q => n6813, QN => n_1474);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n3504, CK => CLK, RN => 
                           RESET, Q => n6814, QN => n_1475);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n3505, CK => CLK, RN => 
                           RESET, Q => n6815, QN => n_1476);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n3506, CK => CLK, RN => 
                           RESET, Q => n6816, QN => n_1477);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n3507, CK => CLK, RN => 
                           RESET, Q => n6817, QN => n_1478);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n3508, CK => CLK, RN => 
                           RESET, Q => n6818, QN => n_1479);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n3509, CK => CLK, RN => 
                           RESET, Q => n6819, QN => n_1480);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n3510, CK => CLK, RN => 
                           RESET, Q => n6820, QN => n_1481);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n3511, CK => CLK, RN => 
                           RESET, Q => n6821, QN => n_1482);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n3512, CK => CLK, RN => 
                           RESET, Q => n6822, QN => n_1483);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n3513, CK => CLK, RN => 
                           RESET, Q => n6823, QN => n_1484);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n3514, CK => CLK, RN => 
                           RESET, Q => n6824, QN => n_1485);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n3515, CK => CLK, RN => 
                           RESET, Q => n6825, QN => n_1486);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n3516, CK => CLK, RN => 
                           RESET, Q => n6826, QN => n_1487);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n3517, CK => CLK, RN => 
                           RESET, Q => n6827, QN => n_1488);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n4093, CK => CLK, RN => 
                           RESET, Q => n7019, QN => n_1489);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n4092, CK => CLK, RN => 
                           RESET, Q => n7018, QN => n_1490);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n4091, CK => CLK, RN => 
                           RESET, Q => n7017, QN => n_1491);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n4090, CK => CLK, RN => 
                           RESET, Q => n7016, QN => n_1492);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n4089, CK => CLK, RN => 
                           RESET, Q => n7015, QN => n_1493);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n4088, CK => CLK, RN => 
                           RESET, Q => n7014, QN => n_1494);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n4087, CK => CLK, RN => 
                           RESET, Q => n7013, QN => n_1495);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n4086, CK => CLK, RN => 
                           RESET, Q => n7012, QN => n_1496);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n4085, CK => CLK, RN => 
                           RESET, Q => n7011, QN => n_1497);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n4084, CK => CLK, RN => 
                           RESET, Q => n7010, QN => n_1498);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n4083, CK => CLK, RN => 
                           RESET, Q => n7009, QN => n_1499);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n4082, CK => CLK, RN => 
                           RESET, Q => n7008, QN => n_1500);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n4081, CK => CLK, RN => 
                           RESET, Q => n7007, QN => n_1501);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n4080, CK => CLK, RN => 
                           RESET, Q => n7006, QN => n_1502);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n4079, CK => CLK, RN => 
                           RESET, Q => n7005, QN => n_1503);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n4078, CK => CLK, RN => 
                           RESET, Q => n7004, QN => n_1504);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n4077, CK => CLK, RN => 
                           RESET, Q => n7003, QN => n_1505);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n4076, CK => CLK, RN => 
                           RESET, Q => n7002, QN => n_1506);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n4075, CK => CLK, RN => 
                           RESET, Q => n7001, QN => n_1507);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n4074, CK => CLK, RN => 
                           RESET, Q => n7000, QN => n_1508);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n4073, CK => CLK, RN => 
                           RESET, Q => n6999, QN => n_1509);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n4072, CK => CLK, RN => 
                           RESET, Q => n6998, QN => n_1510);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n4071, CK => CLK, RN => 
                           RESET, Q => n6997, QN => n_1511);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n4070, CK => CLK, RN => 
                           RESET, Q => n6996, QN => n_1512);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n4069, CK => CLK, RN => 
                           RESET, Q => n6995, QN => n_1513);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n4068, CK => CLK, RN => 
                           RESET, Q => n6994, QN => n_1514);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n4067, CK => CLK, RN => 
                           RESET, Q => n6993, QN => n_1515);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n4066, CK => CLK, RN => 
                           RESET, Q => n6992, QN => n_1516);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n4065, CK => CLK, RN => 
                           RESET, Q => n6991, QN => n_1517);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n4064, CK => CLK, RN => 
                           RESET, Q => n6990, QN => n_1518);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n4063, CK => CLK, RN => 
                           RESET, Q => n6989, QN => n_1519);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n4062, CK => CLK, RN => 
                           RESET, Q => n6988, QN => n_1520);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n4061, CK => CLK, RN => 
                           RESET, Q => n2382, QN => n_1521);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n4060, CK => CLK, RN => 
                           RESET, Q => n2379, QN => n_1522);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n4059, CK => CLK, RN => 
                           RESET, Q => n2376, QN => n_1523);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n4058, CK => CLK, RN => 
                           RESET, Q => n2373, QN => n_1524);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n4057, CK => CLK, RN => 
                           RESET, Q => n2370, QN => n_1525);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n4056, CK => CLK, RN => 
                           RESET, Q => n2367, QN => n_1526);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n4055, CK => CLK, RN => 
                           RESET, Q => n2364, QN => n_1527);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n4054, CK => CLK, RN => 
                           RESET, Q => n2361, QN => n_1528);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n4053, CK => CLK, RN => 
                           RESET, Q => n2358, QN => n_1529);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n4052, CK => CLK, RN => 
                           RESET, Q => n2355, QN => n_1530);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n4051, CK => CLK, RN => 
                           RESET, Q => n2352, QN => n_1531);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n4050, CK => CLK, RN => 
                           RESET, Q => n6763, QN => n_1532);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n4049, CK => CLK, RN => 
                           RESET, Q => n6762, QN => n_1533);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n4048, CK => CLK, RN => 
                           RESET, Q => n6761, QN => n_1534);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n4047, CK => CLK, RN => 
                           RESET, Q => n6760, QN => n_1535);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n4046, CK => CLK, RN => 
                           RESET, Q => n6759, QN => n_1536);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n4045, CK => CLK, RN => 
                           RESET, Q => n6758, QN => n_1537);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n4044, CK => CLK, RN => 
                           RESET, Q => n6757, QN => n_1538);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n4043, CK => CLK, RN => 
                           RESET, Q => n6756, QN => n_1539);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n4042, CK => CLK, RN => 
                           RESET, Q => n6755, QN => n_1540);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n4041, CK => CLK, RN => 
                           RESET, Q => n6754, QN => n_1541);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n4040, CK => CLK, RN => 
                           RESET, Q => n6753, QN => n_1542);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n4039, CK => CLK, RN => 
                           RESET, Q => n6752, QN => n_1543);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n4038, CK => CLK, RN => 
                           RESET, Q => n6751, QN => n_1544);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n4037, CK => CLK, RN => 
                           RESET, Q => n6750, QN => n_1545);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n4036, CK => CLK, RN => 
                           RESET, Q => n6749, QN => n_1546);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n4035, CK => CLK, RN => 
                           RESET, Q => n6748, QN => n_1547);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n4034, CK => CLK, RN => 
                           RESET, Q => n6747, QN => n_1548);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n4033, CK => CLK, RN => 
                           RESET, Q => n6746, QN => n_1549);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n4032, CK => CLK, RN => 
                           RESET, Q => n6745, QN => n_1550);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n4031, CK => CLK, RN => 
                           RESET, Q => n6744, QN => n_1551);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n4030, CK => CLK, RN => 
                           RESET, Q => n6743, QN => n_1552);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n3518, CK => CLK, RN => 
                           RESET, Q => n704, QN => n_1553);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n3519, CK => CLK, RN => 
                           RESET, Q => n703, QN => n_1554);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n3520, CK => CLK, RN => 
                           RESET, Q => n702, QN => n_1555);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n3521, CK => CLK, RN => 
                           RESET, Q => n701, QN => n_1556);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n3522, CK => CLK, RN => 
                           RESET, Q => n700, QN => n_1557);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n3523, CK => CLK, RN => 
                           RESET, Q => n699, QN => n_1558);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n3524, CK => CLK, RN => 
                           RESET, Q => n698, QN => n_1559);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n3525, CK => CLK, RN => 
                           RESET, Q => n697, QN => n_1560);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n3526, CK => CLK, RN => 
                           RESET, Q => n696, QN => n_1561);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n3527, CK => CLK, RN => 
                           RESET, Q => n695, QN => n_1562);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n3528, CK => CLK, RN => 
                           RESET, Q => n694, QN => n_1563);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n3529, CK => CLK, RN => 
                           RESET, Q => n693, QN => n_1564);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n3530, CK => CLK, RN => 
                           RESET, Q => n692, QN => n_1565);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n3531, CK => CLK, RN => 
                           RESET, Q => n691, QN => n_1566);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n3532, CK => CLK, RN => 
                           RESET, Q => n690, QN => n_1567);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n3533, CK => CLK, RN => 
                           RESET, Q => n689, QN => n_1568);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n3534, CK => CLK, RN => 
                           RESET, Q => n688, QN => n_1569);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n3535, CK => CLK, RN => 
                           RESET, Q => n687, QN => n_1570);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n3536, CK => CLK, RN => 
                           RESET, Q => n686, QN => n_1571);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n3537, CK => CLK, RN => 
                           RESET, Q => n685, QN => n_1572);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n3538, CK => CLK, RN => 
                           RESET, Q => n684, QN => n_1573);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n3539, CK => CLK, RN => 
                           RESET, Q => n683, QN => n_1574);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n3540, CK => CLK, RN => 
                           RESET, Q => n682, QN => n_1575);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n3541, CK => CLK, RN => 
                           RESET, Q => n681, QN => n_1576);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n3542, CK => CLK, RN => 
                           RESET, Q => n680, QN => n_1577);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n3543, CK => CLK, RN => 
                           RESET, Q => n679, QN => n_1578);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n3544, CK => CLK, RN => 
                           RESET, Q => n678, QN => n_1579);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n3545, CK => CLK, RN => 
                           RESET, Q => n677, QN => n_1580);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n3546, CK => CLK, RN => 
                           RESET, Q => n676, QN => n_1581);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n3547, CK => CLK, RN => 
                           RESET, Q => n675, QN => n_1582);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n3548, CK => CLK, RN => 
                           RESET, Q => n674, QN => n_1583);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n3549, CK => CLK, RN => 
                           RESET, Q => n673, QN => n_1584);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n3550, CK => CLK, RN => 
                           RESET, Q => n6604, QN => n_1585);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n3551, CK => CLK, RN => 
                           RESET, Q => n6605, QN => n_1586);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n3552, CK => CLK, RN => 
                           RESET, Q => n6606, QN => n_1587);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n3553, CK => CLK, RN => 
                           RESET, Q => n6607, QN => n_1588);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n3554, CK => CLK, RN => 
                           RESET, Q => n6608, QN => n_1589);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n3555, CK => CLK, RN => 
                           RESET, Q => n6609, QN => n_1590);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n3556, CK => CLK, RN => 
                           RESET, Q => n6610, QN => n_1591);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n3557, CK => CLK, RN => 
                           RESET, Q => n6611, QN => n_1592);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n3558, CK => CLK, RN => 
                           RESET, Q => n6612, QN => n_1593);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n3559, CK => CLK, RN => 
                           RESET, Q => n6613, QN => n_1594);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n3560, CK => CLK, RN => 
                           RESET, Q => n6614, QN => n_1595);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n3561, CK => CLK, RN => 
                           RESET, Q => n6615, QN => n_1596);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n3562, CK => CLK, RN => 
                           RESET, Q => n6616, QN => n_1597);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n3563, CK => CLK, RN => 
                           RESET, Q => n6617, QN => n_1598);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n3564, CK => CLK, RN => 
                           RESET, Q => n6618, QN => n_1599);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n3565, CK => CLK, RN => 
                           RESET, Q => n6619, QN => n_1600);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n3566, CK => CLK, RN => 
                           RESET, Q => n6620, QN => n_1601);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n3567, CK => CLK, RN => 
                           RESET, Q => n6621, QN => n_1602);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n3568, CK => CLK, RN => 
                           RESET, Q => n6622, QN => n_1603);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n3569, CK => CLK, RN => 
                           RESET, Q => n6623, QN => n_1604);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n3570, CK => CLK, RN => 
                           RESET, Q => n6624, QN => n_1605);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n3571, CK => CLK, RN => 
                           RESET, Q => n6625, QN => n_1606);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n3572, CK => CLK, RN => 
                           RESET, Q => n6626, QN => n_1607);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n3573, CK => CLK, RN => 
                           RESET, Q => n6627, QN => n_1608);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n3574, CK => CLK, RN => 
                           RESET, Q => n6628, QN => n_1609);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n3575, CK => CLK, RN => 
                           RESET, Q => n6629, QN => n_1610);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n3576, CK => CLK, RN => 
                           RESET, Q => n6630, QN => n_1611);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n3577, CK => CLK, RN => 
                           RESET, Q => n6631, QN => n_1612);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n3578, CK => CLK, RN => 
                           RESET, Q => n6632, QN => n_1613);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n3579, CK => CLK, RN => 
                           RESET, Q => n6633, QN => n_1614);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n3580, CK => CLK, RN => 
                           RESET, Q => n6634, QN => n_1615);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n3581, CK => CLK, RN => 
                           RESET, Q => n6635, QN => n_1616);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n4029, CK => CLK, RN => 
                           RESET, Q => n6707, QN => n_1617);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n4028, CK => CLK, RN => 
                           RESET, Q => n6706, QN => n_1618);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n4027, CK => CLK, RN => 
                           RESET, Q => n6705, QN => n_1619);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n4026, CK => CLK, RN => 
                           RESET, Q => n6704, QN => n_1620);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n4025, CK => CLK, RN => 
                           RESET, Q => n6703, QN => n_1621);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n4024, CK => CLK, RN => 
                           RESET, Q => n6702, QN => n_1622);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n4023, CK => CLK, RN => 
                           RESET, Q => n6701, QN => n_1623);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n4022, CK => CLK, RN => 
                           RESET, Q => n6700, QN => n_1624);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n4021, CK => CLK, RN => 
                           RESET, Q => n6699, QN => n_1625);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n4020, CK => CLK, RN => 
                           RESET, Q => n6698, QN => n_1626);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n4019, CK => CLK, RN => 
                           RESET, Q => n6697, QN => n_1627);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n4018, CK => CLK, RN => 
                           RESET, Q => n6696, QN => n_1628);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n4017, CK => CLK, RN => 
                           RESET, Q => n6695, QN => n_1629);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n4016, CK => CLK, RN => 
                           RESET, Q => n6694, QN => n_1630);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n4015, CK => CLK, RN => 
                           RESET, Q => n6693, QN => n_1631);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n4014, CK => CLK, RN => 
                           RESET, Q => n6692, QN => n_1632);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n4013, CK => CLK, RN => 
                           RESET, Q => n6691, QN => n_1633);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n4012, CK => CLK, RN => 
                           RESET, Q => n6690, QN => n_1634);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n4011, CK => CLK, RN => 
                           RESET, Q => n6689, QN => n_1635);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n4010, CK => CLK, RN => 
                           RESET, Q => n6688, QN => n_1636);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n4009, CK => CLK, RN => 
                           RESET, Q => n6687, QN => n_1637);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n4008, CK => CLK, RN => 
                           RESET, Q => n6686, QN => n_1638);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n4007, CK => CLK, RN => 
                           RESET, Q => n6685, QN => n_1639);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n4006, CK => CLK, RN => 
                           RESET, Q => n6684, QN => n_1640);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n4005, CK => CLK, RN => 
                           RESET, Q => n6683, QN => n_1641);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n4004, CK => CLK, RN => 
                           RESET, Q => n6682, QN => n_1642);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n4003, CK => CLK, RN => 
                           RESET, Q => n6681, QN => n_1643);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n4002, CK => CLK, RN => 
                           RESET, Q => n6680, QN => n_1644);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n4001, CK => CLK, RN => 
                           RESET, Q => n6679, QN => n_1645);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n4000, CK => CLK, RN => 
                           RESET, Q => n6678, QN => n_1646);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n3999, CK => CLK, RN => 
                           RESET, Q => n6677, QN => n_1647);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n3998, CK => CLK, RN => 
                           RESET, Q => n6676, QN => n_1648);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n3790, CK => CLK, RN => 
                           RESET, Q => n6987, QN => n_1649);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n3789, CK => CLK, RN => 
                           RESET, Q => n6986, QN => n_1650);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n3788, CK => CLK, RN => 
                           RESET, Q => n6985, QN => n_1651);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n3787, CK => CLK, RN => 
                           RESET, Q => n6984, QN => n_1652);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n3786, CK => CLK, RN => 
                           RESET, Q => n6983, QN => n_1653);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n3785, CK => CLK, RN => 
                           RESET, Q => n6982, QN => n_1654);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n3784, CK => CLK, RN => 
                           RESET, Q => n6981, QN => n_1655);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n3783, CK => CLK, RN => 
                           RESET, Q => n6980, QN => n_1656);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n3782, CK => CLK, RN => 
                           RESET, Q => n6979, QN => n_1657);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n3781, CK => CLK, RN => 
                           RESET, Q => n6978, QN => n_1658);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n3780, CK => CLK, RN => 
                           RESET, Q => n6977, QN => n_1659);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n3779, CK => CLK, RN => 
                           RESET, Q => n6976, QN => n_1660);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n3778, CK => CLK, RN => 
                           RESET, Q => n6975, QN => n_1661);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n3777, CK => CLK, RN => 
                           RESET, Q => n6974, QN => n_1662);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n3776, CK => CLK, RN => 
                           RESET, Q => n6973, QN => n_1663);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n3775, CK => CLK, RN => 
                           RESET, Q => n6972, QN => n_1664);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n3774, CK => CLK, RN => 
                           RESET, Q => n6971, QN => n_1665);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           RESET, Q => n6904, QN => n_1666);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           RESET, Q => n6901, QN => n_1667);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           RESET, Q => n6898, QN => n_1668);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           RESET, Q => n6895, QN => n_1669);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           RESET, Q => n6892, QN => n_1670);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           RESET, Q => n6889, QN => n_1671);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           RESET, Q => n6886, QN => n_1672);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           RESET, Q => n6883, QN => n_1673);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           RESET, Q => n6880, QN => n_1674);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           RESET, Q => n6877, QN => n_1675);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           RESET, Q => n6874, QN => n_1676);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           RESET, Q => n6871, QN => n_1677);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           RESET, Q => n6868, QN => n_1678);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           RESET, Q => n6865, QN => n_1679);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           RESET, Q => n6862, QN => n_1680);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n3582, CK => CLK, RN => 
                           RESET, Q => n736, QN => n_1681);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n3583, CK => CLK, RN => 
                           RESET, Q => n735, QN => n_1682);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n3584, CK => CLK, RN => 
                           RESET, Q => n734, QN => n_1683);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n3585, CK => CLK, RN => 
                           RESET, Q => n733, QN => n_1684);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n3586, CK => CLK, RN => 
                           RESET, Q => n732, QN => n_1685);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n3587, CK => CLK, RN => 
                           RESET, Q => n731, QN => n_1686);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n3588, CK => CLK, RN => 
                           RESET, Q => n730, QN => n_1687);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n3589, CK => CLK, RN => 
                           RESET, Q => n729, QN => n_1688);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n3590, CK => CLK, RN => 
                           RESET, Q => n728, QN => n_1689);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n3591, CK => CLK, RN => 
                           RESET, Q => n727, QN => n_1690);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n3592, CK => CLK, RN => 
                           RESET, Q => n726, QN => n_1691);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n3593, CK => CLK, RN => 
                           RESET, Q => n725, QN => n_1692);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n3594, CK => CLK, RN => 
                           RESET, Q => n724, QN => n_1693);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n3595, CK => CLK, RN => 
                           RESET, Q => n723, QN => n_1694);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n3596, CK => CLK, RN => 
                           RESET, Q => n722, QN => n_1695);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n3597, CK => CLK, RN => 
                           RESET, Q => n721, QN => n_1696);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n3598, CK => CLK, RN => 
                           RESET, Q => n720, QN => n_1697);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n3599, CK => CLK, RN => 
                           RESET, Q => n719, QN => n_1698);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n3600, CK => CLK, RN => 
                           RESET, Q => n718, QN => n_1699);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n3601, CK => CLK, RN => 
                           RESET, Q => n717, QN => n_1700);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n3602, CK => CLK, RN => 
                           RESET, Q => n716, QN => n_1701);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n3603, CK => CLK, RN => 
                           RESET, Q => n715, QN => n_1702);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n3604, CK => CLK, RN => 
                           RESET, Q => n714, QN => n_1703);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n3605, CK => CLK, RN => 
                           RESET, Q => n713, QN => n_1704);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n3606, CK => CLK, RN => 
                           RESET, Q => n712, QN => n_1705);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n3607, CK => CLK, RN => 
                           RESET, Q => n711, QN => n_1706);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n3608, CK => CLK, RN => 
                           RESET, Q => n710, QN => n_1707);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n3609, CK => CLK, RN => 
                           RESET, Q => n709, QN => n_1708);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n3610, CK => CLK, RN => 
                           RESET, Q => n708, QN => n_1709);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n3611, CK => CLK, RN => 
                           RESET, Q => n707, QN => n_1710);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n3612, CK => CLK, RN => 
                           RESET, Q => n706, QN => n_1711);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n3613, CK => CLK, RN => 
                           RESET, Q => n705, QN => n_1712);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n3614, CK => CLK, RN => 
                           RESET, Q => n544, QN => n_1713);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n3615, CK => CLK, RN => 
                           RESET, Q => n543, QN => n_1714);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n3616, CK => CLK, RN => 
                           RESET, Q => n542, QN => n_1715);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n3617, CK => CLK, RN => 
                           RESET, Q => n541, QN => n_1716);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n3618, CK => CLK, RN => 
                           RESET, Q => n540, QN => n_1717);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n3619, CK => CLK, RN => 
                           RESET, Q => n539, QN => n_1718);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n3620, CK => CLK, RN => 
                           RESET, Q => n538, QN => n_1719);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n3621, CK => CLK, RN => 
                           RESET, Q => n537, QN => n_1720);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n3622, CK => CLK, RN => 
                           RESET, Q => n536, QN => n_1721);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n3623, CK => CLK, RN => 
                           RESET, Q => n535, QN => n_1722);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n3624, CK => CLK, RN => 
                           RESET, Q => n534, QN => n_1723);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n3625, CK => CLK, RN => 
                           RESET, Q => n533, QN => n_1724);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n3626, CK => CLK, RN => 
                           RESET, Q => n532, QN => n_1725);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n3627, CK => CLK, RN => 
                           RESET, Q => n531, QN => n_1726);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n3628, CK => CLK, RN => 
                           RESET, Q => n530, QN => n_1727);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n3629, CK => CLK, RN => 
                           RESET, Q => n529, QN => n_1728);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n3630, CK => CLK, RN => 
                           RESET, Q => n528, QN => n_1729);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n3631, CK => CLK, RN => 
                           RESET, Q => n527, QN => n_1730);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n3632, CK => CLK, RN => 
                           RESET, Q => n526, QN => n_1731);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n3633, CK => CLK, RN => 
                           RESET, Q => n525, QN => n_1732);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n3634, CK => CLK, RN => 
                           RESET, Q => n524, QN => n_1733);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n3635, CK => CLK, RN => 
                           RESET, Q => n523, QN => n_1734);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n3636, CK => CLK, RN => 
                           RESET, Q => n522, QN => n_1735);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n3637, CK => CLK, RN => 
                           RESET, Q => n521, QN => n_1736);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n3638, CK => CLK, RN => 
                           RESET, Q => n520, QN => n_1737);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n3639, CK => CLK, RN => 
                           RESET, Q => n519, QN => n_1738);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n3640, CK => CLK, RN => 
                           RESET, Q => n518, QN => n_1739);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n3641, CK => CLK, RN => 
                           RESET, Q => n517, QN => n_1740);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n3642, CK => CLK, RN => 
                           RESET, Q => n516, QN => n_1741);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n3643, CK => CLK, RN => 
                           RESET, Q => n515, QN => n_1742);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n3644, CK => CLK, RN => 
                           RESET, Q => n514, QN => n_1743);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n3645, CK => CLK, RN => 
                           RESET, Q => n513, QN => n_1744);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n3886, CK => CLK, RN => 
                           RESET, Q => n6859, QN => n_1745);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n3885, CK => CLK, RN => 
                           RESET, Q => n6858, QN => n_1746);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n3884, CK => CLK, RN => 
                           RESET, Q => n6857, QN => n_1747);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n3883, CK => CLK, RN => 
                           RESET, Q => n6856, QN => n_1748);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n3882, CK => CLK, RN => 
                           RESET, Q => n6855, QN => n_1749);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n3881, CK => CLK, RN => 
                           RESET, Q => n6854, QN => n_1750);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n3880, CK => CLK, RN => 
                           RESET, Q => n6853, QN => n_1751);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n3879, CK => CLK, RN => 
                           RESET, Q => n6852, QN => n_1752);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n3878, CK => CLK, RN => 
                           RESET, Q => n6851, QN => n_1753);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n3877, CK => CLK, RN => 
                           RESET, Q => n6850, QN => n_1754);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n3876, CK => CLK, RN => 
                           RESET, Q => n6849, QN => n_1755);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n3875, CK => CLK, RN => 
                           RESET, Q => n6848, QN => n_1756);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n3874, CK => CLK, RN => 
                           RESET, Q => n6847, QN => n_1757);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n3873, CK => CLK, RN => 
                           RESET, Q => n6846, QN => n_1758);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n3872, CK => CLK, RN => 
                           RESET, Q => n6845, QN => n_1759);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n3871, CK => CLK, RN => 
                           RESET, Q => n6844, QN => n_1760);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n3870, CK => CLK, RN => 
                           RESET, Q => n6843, QN => n_1761);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n3805, CK => CLK, RN => 
                           RESET, Q => n6842, QN => n_1762);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n3804, CK => CLK, RN => 
                           RESET, Q => n6841, QN => n_1763);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n3803, CK => CLK, RN => 
                           RESET, Q => n6840, QN => n_1764);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n3802, CK => CLK, RN => 
                           RESET, Q => n6839, QN => n_1765);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n3801, CK => CLK, RN => 
                           RESET, Q => n6838, QN => n_1766);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n3800, CK => CLK, RN => 
                           RESET, Q => n6837, QN => n_1767);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n3799, CK => CLK, RN => 
                           RESET, Q => n6836, QN => n_1768);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n3798, CK => CLK, RN => 
                           RESET, Q => n6835, QN => n_1769);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n3797, CK => CLK, RN => 
                           RESET, Q => n6834, QN => n_1770);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n3796, CK => CLK, RN => 
                           RESET, Q => n6833, QN => n_1771);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n3795, CK => CLK, RN => 
                           RESET, Q => n6832, QN => n_1772);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n3794, CK => CLK, RN => 
                           RESET, Q => n6831, QN => n_1773);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n3793, CK => CLK, RN => 
                           RESET, Q => n6830, QN => n_1774);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n3792, CK => CLK, RN => 
                           RESET, Q => n6829, QN => n_1775);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n3791, CK => CLK, RN => 
                           RESET, Q => n6828, QN => n_1776);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n3918, CK => CLK, RN => 
                           RESET, Q => n7115, QN => n1423);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n3917, CK => CLK, RN => 
                           RESET, Q => n7114, QN => n1424);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n3916, CK => CLK, RN => 
                           RESET, Q => n7113, QN => n1425);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n3915, CK => CLK, RN => 
                           RESET, Q => n7112, QN => n1426);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n3914, CK => CLK, RN => 
                           RESET, Q => n7111, QN => n1427);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n3913, CK => CLK, RN => 
                           RESET, Q => n7110, QN => n1428);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n3912, CK => CLK, RN => 
                           RESET, Q => n7109, QN => n1429);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n3911, CK => CLK, RN => 
                           RESET, Q => n7108, QN => n1430);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n3910, CK => CLK, RN => 
                           RESET, Q => n7107, QN => n1431);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n3909, CK => CLK, RN => 
                           RESET, Q => n7106, QN => n1432);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n3908, CK => CLK, RN => 
                           RESET, Q => n7105, QN => n1433);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n3907, CK => CLK, RN => 
                           RESET, Q => n7104, QN => n1434);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n3906, CK => CLK, RN => 
                           RESET, Q => n7103, QN => n1435);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n3905, CK => CLK, RN => 
                           RESET, Q => n7102, QN => n1436);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n3904, CK => CLK, RN => 
                           RESET, Q => n7101, QN => n1437);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n3903, CK => CLK, RN => 
                           RESET, Q => n7100, QN => n1438);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n3902, CK => CLK, RN => 
                           RESET, Q => n7099, QN => n1439);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n3901, CK => CLK, RN => 
                           RESET, Q => n7098, QN => n1440);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n3900, CK => CLK, RN => 
                           RESET, Q => n7097, QN => n1441);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n3899, CK => CLK, RN => 
                           RESET, Q => n7096, QN => n1442);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n3898, CK => CLK, RN => 
                           RESET, Q => n7095, QN => n1443);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n3897, CK => CLK, RN => 
                           RESET, Q => n7094, QN => n1444);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n3896, CK => CLK, RN => 
                           RESET, Q => n7093, QN => n1445);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n3895, CK => CLK, RN => 
                           RESET, Q => n7092, QN => n1446);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n3894, CK => CLK, RN => 
                           RESET, Q => n7091, QN => n1447);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n3893, CK => CLK, RN => 
                           RESET, Q => n7090, QN => n1448);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n3892, CK => CLK, RN => 
                           RESET, Q => n7089, QN => n1449);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n3891, CK => CLK, RN => 
                           RESET, Q => n7088, QN => n1450);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n3890, CK => CLK, RN => 
                           RESET, Q => n7087, QN => n1451);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n3889, CK => CLK, RN => 
                           RESET, Q => n7086, QN => n1452);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n3888, CK => CLK, RN => 
                           RESET, Q => n7085, QN => n1453);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n3887, CK => CLK, RN => 
                           RESET, Q => n7084, QN => n1454);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           RESET, Q => n6938, QN => n_1777);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           RESET, Q => n6936, QN => n_1778);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           RESET, Q => n6934, QN => n_1779);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           RESET, Q => n6932, QN => n_1780);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           RESET, Q => n6930, QN => n_1781);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           RESET, Q => n6928, QN => n_1782);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           RESET, Q => n6926, QN => n_1783);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           RESET, Q => n6924, QN => n_1784);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           RESET, Q => n6922, QN => n_1785);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           RESET, Q => n6920, QN => n_1786);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           RESET, Q => n6918, QN => n_1787);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           RESET, Q => n6916, QN => n_1788);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           RESET, Q => n6914, QN => n_1789);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           RESET, Q => n6912, QN => n_1790);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           RESET, Q => n6910, QN => n_1791);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           RESET, Q => n6908, QN => n_1792);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           RESET, Q => n6906, QN => n_1793);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           RESET, Q => n6903, QN => n_1794);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           RESET, Q => n6900, QN => n_1795);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           RESET, Q => n6897, QN => n_1796);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           RESET, Q => n6894, QN => n_1797);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           RESET, Q => n6891, QN => n_1798);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           RESET, Q => n6888, QN => n_1799);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           RESET, Q => n6885, QN => n_1800);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           RESET, Q => n6882, QN => n_1801);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           RESET, Q => n6879, QN => n_1802);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           RESET, Q => n6876, QN => n_1803);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           RESET, Q => n6873, QN => n_1804);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           RESET, Q => n6870, QN => n_1805);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           RESET, Q => n6867, QN => n_1806);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           RESET, Q => n6864, QN => n_1807);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           RESET, Q => n6861, QN => n_1808);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n3869, CK => CLK, RN => 
                           RESET, Q => n2830, QN => n_1809);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n3868, CK => CLK, RN => 
                           RESET, Q => n2829, QN => n_1810);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n3867, CK => CLK, RN => 
                           RESET, Q => n2828, QN => n_1811);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n3866, CK => CLK, RN => 
                           RESET, Q => n2827, QN => n_1812);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n3865, CK => CLK, RN => 
                           RESET, Q => n2826, QN => n_1813);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n3864, CK => CLK, RN => 
                           RESET, Q => n2825, QN => n_1814);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n3863, CK => CLK, RN => 
                           RESET, Q => n2824, QN => n_1815);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n3862, CK => CLK, RN => 
                           RESET, Q => n2823, QN => n_1816);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n3861, CK => CLK, RN => 
                           RESET, Q => n2822, QN => n_1817);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n3860, CK => CLK, RN => 
                           RESET, Q => n2821, QN => n_1818);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n3859, CK => CLK, RN => 
                           RESET, Q => n2820, QN => n_1819);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n3858, CK => CLK, RN => 
                           RESET, Q => n2819, QN => n_1820);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n3857, CK => CLK, RN => 
                           RESET, Q => n2818, QN => n_1821);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n3856, CK => CLK, RN => 
                           RESET, Q => n2817, QN => n_1822);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n3855, CK => CLK, RN => 
                           RESET, Q => n2816, QN => n_1823);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n3854, CK => CLK, RN => 
                           RESET, Q => n2815, QN => n_1824);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n3853, CK => CLK, RN => 
                           RESET, Q => n2814, QN => n_1825);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n3852, CK => CLK, RN => 
                           RESET, Q => n2813, QN => n_1826);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n3851, CK => CLK, RN => 
                           RESET, Q => n2812, QN => n_1827);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n3850, CK => CLK, RN => 
                           RESET, Q => n2811, QN => n_1828);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n3849, CK => CLK, RN => 
                           RESET, Q => n2810, QN => n_1829);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n3848, CK => CLK, RN => 
                           RESET, Q => n2809, QN => n_1830);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n3847, CK => CLK, RN => 
                           RESET, Q => n2808, QN => n_1831);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n3846, CK => CLK, RN => 
                           RESET, Q => n2807, QN => n_1832);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n3845, CK => CLK, RN => 
                           RESET, Q => n6675, QN => n_1833);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n3844, CK => CLK, RN => 
                           RESET, Q => n6674, QN => n_1834);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n3843, CK => CLK, RN => 
                           RESET, Q => n6673, QN => n_1835);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n3842, CK => CLK, RN => 
                           RESET, Q => n6672, QN => n_1836);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n3841, CK => CLK, RN => 
                           RESET, Q => n6671, QN => n_1837);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n3840, CK => CLK, RN => 
                           RESET, Q => n6670, QN => n_1838);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n3839, CK => CLK, RN => 
                           RESET, Q => n6669, QN => n_1839);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n3838, CK => CLK, RN => 
                           RESET, Q => n6668, QN => n_1840);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n3646, CK => CLK, RN => 
                           RESET, Q => n512, QN => n_1841);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n3647, CK => CLK, RN => 
                           RESET, Q => n511, QN => n_1842);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n3648, CK => CLK, RN => 
                           RESET, Q => n510, QN => n_1843);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n3649, CK => CLK, RN => 
                           RESET, Q => n509, QN => n_1844);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n3650, CK => CLK, RN => 
                           RESET, Q => n508, QN => n_1845);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n3651, CK => CLK, RN => 
                           RESET, Q => n507, QN => n_1846);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n3652, CK => CLK, RN => 
                           RESET, Q => n506, QN => n_1847);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n3653, CK => CLK, RN => 
                           RESET, Q => n505, QN => n_1848);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n3654, CK => CLK, RN => 
                           RESET, Q => n504, QN => n_1849);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n3655, CK => CLK, RN => 
                           RESET, Q => n503, QN => n_1850);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n3656, CK => CLK, RN => 
                           RESET, Q => n502, QN => n_1851);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n3657, CK => CLK, RN => 
                           RESET, Q => n501, QN => n_1852);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n3658, CK => CLK, RN => 
                           RESET, Q => n500, QN => n_1853);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n3659, CK => CLK, RN => 
                           RESET, Q => n499, QN => n_1854);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n3660, CK => CLK, RN => 
                           RESET, Q => n498, QN => n_1855);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n3661, CK => CLK, RN => 
                           RESET, Q => n497, QN => n_1856);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n3662, CK => CLK, RN => 
                           RESET, Q => n496, QN => n_1857);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n3663, CK => CLK, RN => 
                           RESET, Q => n495, QN => n_1858);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n3664, CK => CLK, RN => 
                           RESET, Q => n494, QN => n_1859);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n3665, CK => CLK, RN => 
                           RESET, Q => n493, QN => n_1860);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n3666, CK => CLK, RN => 
                           RESET, Q => n492, QN => n_1861);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n3667, CK => CLK, RN => 
                           RESET, Q => n491, QN => n_1862);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n3668, CK => CLK, RN => 
                           RESET, Q => n490, QN => n_1863);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n3669, CK => CLK, RN => 
                           RESET, Q => n489, QN => n_1864);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n3670, CK => CLK, RN => 
                           RESET, Q => n488, QN => n_1865);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n3671, CK => CLK, RN => 
                           RESET, Q => n487, QN => n_1866);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n3672, CK => CLK, RN => 
                           RESET, Q => n486, QN => n_1867);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n3673, CK => CLK, RN => 
                           RESET, Q => n485, QN => n_1868);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n3674, CK => CLK, RN => 
                           RESET, Q => n484, QN => n_1869);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n3675, CK => CLK, RN => 
                           RESET, Q => n483, QN => n_1870);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n3676, CK => CLK, RN => 
                           RESET, Q => n482, QN => n_1871);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n3677, CK => CLK, RN => 
                           RESET, Q => n481, QN => n_1872);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n3678, CK => CLK, RN => 
                           RESET, Q => n672, QN => n_1873);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n3679, CK => CLK, RN => 
                           RESET, Q => n671, QN => n_1874);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n3680, CK => CLK, RN => 
                           RESET, Q => n670, QN => n_1875);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n3681, CK => CLK, RN => 
                           RESET, Q => n669, QN => n_1876);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n3682, CK => CLK, RN => 
                           RESET, Q => n668, QN => n_1877);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n3683, CK => CLK, RN => 
                           RESET, Q => n667, QN => n_1878);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n3684, CK => CLK, RN => 
                           RESET, Q => n666, QN => n_1879);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n3685, CK => CLK, RN => 
                           RESET, Q => n665, QN => n_1880);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n3686, CK => CLK, RN => 
                           RESET, Q => n664, QN => n_1881);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n3687, CK => CLK, RN => 
                           RESET, Q => n663, QN => n_1882);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n3688, CK => CLK, RN => 
                           RESET, Q => n662, QN => n_1883);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n3689, CK => CLK, RN => 
                           RESET, Q => n661, QN => n_1884);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n3690, CK => CLK, RN => 
                           RESET, Q => n660, QN => n_1885);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n3691, CK => CLK, RN => 
                           RESET, Q => n659, QN => n_1886);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n3692, CK => CLK, RN => 
                           RESET, Q => n658, QN => n_1887);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n3693, CK => CLK, RN => 
                           RESET, Q => n657, QN => n_1888);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n3694, CK => CLK, RN => 
                           RESET, Q => n656, QN => n_1889);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n3695, CK => CLK, RN => 
                           RESET, Q => n655, QN => n_1890);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n3696, CK => CLK, RN => 
                           RESET, Q => n654, QN => n_1891);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n3697, CK => CLK, RN => 
                           RESET, Q => n653, QN => n_1892);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n3698, CK => CLK, RN => 
                           RESET, Q => n652, QN => n_1893);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n3699, CK => CLK, RN => 
                           RESET, Q => n651, QN => n_1894);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n3700, CK => CLK, RN => 
                           RESET, Q => n650, QN => n_1895);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n3701, CK => CLK, RN => 
                           RESET, Q => n649, QN => n_1896);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n3702, CK => CLK, RN => 
                           RESET, Q => n648, QN => n_1897);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n3703, CK => CLK, RN => 
                           RESET, Q => n647, QN => n_1898);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n3704, CK => CLK, RN => 
                           RESET, Q => n646, QN => n_1899);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n3705, CK => CLK, RN => 
                           RESET, Q => n645, QN => n_1900);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n3706, CK => CLK, RN => 
                           RESET, Q => n644, QN => n_1901);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n3707, CK => CLK, RN => 
                           RESET, Q => n643, QN => n_1902);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n3708, CK => CLK, RN => 
                           RESET, Q => n642, QN => n_1903);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n3709, CK => CLK, RN => 
                           RESET, Q => n641, QN => n_1904);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n3837, CK => CLK, RN => 
                           RESET, Q => n6742, QN => n_1905);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n3836, CK => CLK, RN => 
                           RESET, Q => n6741, QN => n_1906);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n3835, CK => CLK, RN => 
                           RESET, Q => n6740, QN => n_1907);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n3834, CK => CLK, RN => 
                           RESET, Q => n6739, QN => n_1908);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n3833, CK => CLK, RN => 
                           RESET, Q => n6738, QN => n_1909);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n3832, CK => CLK, RN => 
                           RESET, Q => n6737, QN => n_1910);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n3831, CK => CLK, RN => 
                           RESET, Q => n6736, QN => n_1911);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n3830, CK => CLK, RN => 
                           RESET, Q => n6735, QN => n_1912);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n3829, CK => CLK, RN => 
                           RESET, Q => n6734, QN => n_1913);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n3828, CK => CLK, RN => 
                           RESET, Q => n6733, QN => n_1914);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n3827, CK => CLK, RN => 
                           RESET, Q => n6732, QN => n_1915);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n3826, CK => CLK, RN => 
                           RESET, Q => n6731, QN => n_1916);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n3825, CK => CLK, RN => 
                           RESET, Q => n6730, QN => n_1917);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n3824, CK => CLK, RN => 
                           RESET, Q => n6729, QN => n_1918);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n3823, CK => CLK, RN => 
                           RESET, Q => n6728, QN => n_1919);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n3822, CK => CLK, RN => 
                           RESET, Q => n6727, QN => n_1920);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n3821, CK => CLK, RN => 
                           RESET, Q => n6726, QN => n_1921);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n3820, CK => CLK, RN => 
                           RESET, Q => n6725, QN => n_1922);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n3819, CK => CLK, RN => 
                           RESET, Q => n6724, QN => n_1923);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n3818, CK => CLK, RN => 
                           RESET, Q => n6723, QN => n_1924);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n3817, CK => CLK, RN => 
                           RESET, Q => n6722, QN => n_1925);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n3816, CK => CLK, RN => 
                           RESET, Q => n6721, QN => n_1926);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n3815, CK => CLK, RN => 
                           RESET, Q => n6720, QN => n_1927);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n3814, CK => CLK, RN => 
                           RESET, Q => n6719, QN => n_1928);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n3813, CK => CLK, RN => 
                           RESET, Q => n6718, QN => n_1929);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n3812, CK => CLK, RN => 
                           RESET, Q => n6717, QN => n_1930);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n3811, CK => CLK, RN => 
                           RESET, Q => n6716, QN => n_1931);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n3810, CK => CLK, RN => 
                           RESET, Q => n6715, QN => n_1932);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n3809, CK => CLK, RN => 
                           RESET, Q => n6714, QN => n_1933);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n3808, CK => CLK, RN => 
                           RESET, Q => n6713, QN => n_1934);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n3807, CK => CLK, RN => 
                           RESET, Q => n6712, QN => n_1935);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n3806, CK => CLK, RN => 
                           RESET, Q => n6711, QN => n_1936);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           RESET, Q => n6937, QN => n_1937);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           RESET, Q => n6935, QN => n_1938);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           RESET, Q => n6933, QN => n_1939);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           RESET, Q => n6931, QN => n_1940);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           RESET, Q => n6929, QN => n_1941);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           RESET, Q => n6927, QN => n_1942);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           RESET, Q => n6925, QN => n_1943);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           RESET, Q => n6923, QN => n_1944);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           RESET, Q => n6921, QN => n_1945);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           RESET, Q => n6919, QN => n_1946);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           RESET, Q => n6917, QN => n_1947);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           RESET, Q => n6915, QN => n_1948);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           RESET, Q => n6913, QN => n_1949);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           RESET, Q => n6911, QN => n_1950);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           RESET, Q => n6909, QN => n_1951);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           RESET, Q => n6907, QN => n_1952);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           RESET, Q => n6905, QN => n_1953);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           RESET, Q => n6902, QN => n_1954);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           RESET, Q => n6899, QN => n_1955);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           RESET, Q => n6896, QN => n_1956);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           RESET, Q => n6893, QN => n_1957);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           RESET, Q => n6890, QN => n_1958);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           RESET, Q => n6887, QN => n_1959);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           RESET, Q => n6884, QN => n_1960);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           RESET, Q => n6881, QN => n_1961);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           RESET, Q => n6878, QN => n_1962);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           RESET, Q => n6875, QN => n_1963);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           RESET, Q => n6872, QN => n_1964);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           RESET, Q => n6869, QN => n_1965);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           RESET, Q => n6866, QN => n_1966);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           RESET, Q => n6863, QN => n_1967);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           RESET, Q => n6860, QN => n_1968);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n3710, CK => CLK, RN => 
                           RESET, Q => n384, QN => n_1969);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n3711, CK => CLK, RN => 
                           RESET, Q => n383, QN => n_1970);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n3712, CK => CLK, RN => 
                           RESET, Q => n382, QN => n_1971);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n3713, CK => CLK, RN => 
                           RESET, Q => n381, QN => n_1972);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n3714, CK => CLK, RN => 
                           RESET, Q => n380, QN => n_1973);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n3715, CK => CLK, RN => 
                           RESET, Q => n379, QN => n_1974);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n3716, CK => CLK, RN => 
                           RESET, Q => n378, QN => n_1975);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n3717, CK => CLK, RN => 
                           RESET, Q => n377, QN => n_1976);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n3718, CK => CLK, RN => 
                           RESET, Q => n376, QN => n_1977);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n3719, CK => CLK, RN => 
                           RESET, Q => n375, QN => n_1978);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n3720, CK => CLK, RN => 
                           RESET, Q => n374, QN => n_1979);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n3721, CK => CLK, RN => 
                           RESET, Q => n373, QN => n_1980);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n3722, CK => CLK, RN => 
                           RESET, Q => n372, QN => n_1981);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n3723, CK => CLK, RN => 
                           RESET, Q => n371, QN => n_1982);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n3724, CK => CLK, RN => 
                           RESET, Q => n370, QN => n_1983);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n3725, CK => CLK, RN => 
                           RESET, Q => n369, QN => n_1984);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n3726, CK => CLK, RN => 
                           RESET, Q => n368, QN => n_1985);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n3727, CK => CLK, RN => 
                           RESET, Q => n367, QN => n_1986);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n3728, CK => CLK, RN => 
                           RESET, Q => n366, QN => n_1987);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n3729, CK => CLK, RN => 
                           RESET, Q => n365, QN => n_1988);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n3730, CK => CLK, RN => 
                           RESET, Q => n364, QN => n_1989);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n3731, CK => CLK, RN => 
                           RESET, Q => n363, QN => n_1990);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n3732, CK => CLK, RN => 
                           RESET, Q => n362, QN => n_1991);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n3733, CK => CLK, RN => 
                           RESET, Q => n361, QN => n_1992);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n3734, CK => CLK, RN => 
                           RESET, Q => n360, QN => n_1993);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n3735, CK => CLK, RN => 
                           RESET, Q => n359, QN => n_1994);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n3736, CK => CLK, RN => 
                           RESET, Q => n358, QN => n_1995);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n3737, CK => CLK, RN => 
                           RESET, Q => n357, QN => n_1996);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n3738, CK => CLK, RN => 
                           RESET, Q => n356, QN => n_1997);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n3739, CK => CLK, RN => 
                           RESET, Q => n355, QN => n_1998);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n3740, CK => CLK, RN => 
                           RESET, Q => n354, QN => n_1999);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n3741, CK => CLK, RN => 
                           RESET, Q => n353, QN => n_2000);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n3742, CK => CLK, RN => 
                           RESET, Q => n352, QN => n_2001);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n3743, CK => CLK, RN => 
                           RESET, Q => n351, QN => n_2002);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n3744, CK => CLK, RN => 
                           RESET, Q => n350, QN => n_2003);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n3745, CK => CLK, RN => 
                           RESET, Q => n349, QN => n_2004);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n3746, CK => CLK, RN => 
                           RESET, Q => n348, QN => n_2005);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n3747, CK => CLK, RN => 
                           RESET, Q => n347, QN => n_2006);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n3748, CK => CLK, RN => 
                           RESET, Q => n346, QN => n_2007);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n3749, CK => CLK, RN => 
                           RESET, Q => n345, QN => n_2008);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n3750, CK => CLK, RN => 
                           RESET, Q => n344, QN => n_2009);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n3751, CK => CLK, RN => 
                           RESET, Q => n343, QN => n_2010);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n3752, CK => CLK, RN => 
                           RESET, Q => n342, QN => n_2011);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n3753, CK => CLK, RN => 
                           RESET, Q => n341, QN => n_2012);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n3754, CK => CLK, RN => 
                           RESET, Q => n340, QN => n_2013);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n3755, CK => CLK, RN => 
                           RESET, Q => n339, QN => n_2014);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n3756, CK => CLK, RN => 
                           RESET, Q => n338, QN => n_2015);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n3757, CK => CLK, RN => 
                           RESET, Q => n337, QN => n_2016);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n3758, CK => CLK, RN => 
                           RESET, Q => n336, QN => n_2017);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n3759, CK => CLK, RN => 
                           RESET, Q => n335, QN => n_2018);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n3760, CK => CLK, RN => 
                           RESET, Q => n334, QN => n_2019);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n3761, CK => CLK, RN => 
                           RESET, Q => n333, QN => n_2020);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n3762, CK => CLK, RN => 
                           RESET, Q => n332, QN => n_2021);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n3763, CK => CLK, RN => 
                           RESET, Q => n331, QN => n_2022);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n3764, CK => CLK, RN => 
                           RESET, Q => n330, QN => n_2023);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n3765, CK => CLK, RN => 
                           RESET, Q => n329, QN => n_2024);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n3766, CK => CLK, RN => 
                           RESET, Q => n328, QN => n_2025);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n3767, CK => CLK, RN => 
                           RESET, Q => n327, QN => n_2026);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n3768, CK => CLK, RN => 
                           RESET, Q => n326, QN => n_2027);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n3769, CK => CLK, RN => 
                           RESET, Q => n325, QN => n_2028);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n3770, CK => CLK, RN => 
                           RESET, Q => n324, QN => n_2029);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n3771, CK => CLK, RN => 
                           RESET, Q => n323, QN => n_2030);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n3772, CK => CLK, RN => 
                           RESET, Q => n322, QN => n_2031);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n3773, CK => CLK, RN => 
                           RESET, Q => n321, QN => n_2032);
   OUT1_reg_31_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => RESET, Q 
                           => OUT1_31_port, QN => n_2033);
   OUT1_reg_30_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => RESET, Q 
                           => OUT1_30_port, QN => n_2034);
   OUT1_reg_29_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => RESET, Q 
                           => OUT1_29_port, QN => n_2035);
   OUT1_reg_28_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => RESET, Q 
                           => OUT1_28_port, QN => n_2036);
   OUT1_reg_27_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => RESET, Q 
                           => OUT1_27_port, QN => n_2037);
   OUT1_reg_26_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => RESET, Q 
                           => OUT1_26_port, QN => n_2038);
   OUT1_reg_25_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => RESET, Q 
                           => OUT1_25_port, QN => n_2039);
   OUT1_reg_24_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => RESET, Q 
                           => OUT1_24_port, QN => n_2040);
   OUT1_reg_23_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => RESET, Q 
                           => OUT1_23_port, QN => n_2041);
   OUT1_reg_22_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => RESET, Q 
                           => OUT1_22_port, QN => n_2042);
   OUT1_reg_21_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => RESET, Q 
                           => OUT1_21_port, QN => n_2043);
   OUT1_reg_20_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => RESET, Q 
                           => OUT1_20_port, QN => n_2044);
   OUT1_reg_19_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => RESET, Q 
                           => OUT1_19_port, QN => n_2045);
   OUT1_reg_18_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => RESET, Q 
                           => OUT1_18_port, QN => n_2046);
   OUT1_reg_17_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => RESET, Q 
                           => OUT1_17_port, QN => n_2047);
   OUT1_reg_16_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => RESET, Q 
                           => OUT1_16_port, QN => n_2048);
   OUT1_reg_15_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => RESET, Q 
                           => OUT1_15_port, QN => n_2049);
   OUT1_reg_14_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => RESET, Q 
                           => OUT1_14_port, QN => n_2050);
   OUT1_reg_13_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => RESET, Q 
                           => OUT1_13_port, QN => n_2051);
   OUT1_reg_12_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => RESET, Q 
                           => OUT1_12_port, QN => n_2052);
   OUT1_reg_11_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => RESET, Q 
                           => OUT1_11_port, QN => n_2053);
   OUT1_reg_10_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => RESET, Q 
                           => OUT1_10_port, QN => n_2054);
   OUT1_reg_9_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => RESET, Q =>
                           OUT1_9_port, QN => n_2055);
   OUT1_reg_8_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => RESET, Q =>
                           OUT1_8_port, QN => n_2056);
   OUT1_reg_7_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => RESET, Q =>
                           OUT1_7_port, QN => n_2057);
   OUT1_reg_6_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => RESET, Q =>
                           OUT1_6_port, QN => n_2058);
   OUT1_reg_5_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => RESET, Q =>
                           OUT1_5_port, QN => n_2059);
   OUT1_reg_4_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => RESET, Q =>
                           OUT1_4_port, QN => n_2060);
   OUT1_reg_3_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => RESET, Q =>
                           OUT1_3_port, QN => n_2061);
   OUT1_reg_2_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => RESET, Q =>
                           OUT1_2_port, QN => n_2062);
   OUT1_reg_1_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => RESET, Q =>
                           OUT1_1_port, QN => n_2063);
   OUT1_reg_0_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => RESET, Q =>
                           OUT1_0_port, QN => n_2064);
   OUT2_reg_31_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => RESET, Q 
                           => OUT2_31_port, QN => n_2065);
   OUT2_reg_30_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => RESET, Q 
                           => OUT2_30_port, QN => n_2066);
   OUT2_reg_29_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => RESET, Q 
                           => OUT2_29_port, QN => n_2067);
   OUT2_reg_28_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => RESET, Q 
                           => OUT2_28_port, QN => n_2068);
   OUT2_reg_27_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => RESET, Q 
                           => OUT2_27_port, QN => n_2069);
   OUT2_reg_26_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => RESET, Q 
                           => OUT2_26_port, QN => n_2070);
   OUT2_reg_25_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => RESET, Q 
                           => OUT2_25_port, QN => n_2071);
   OUT2_reg_24_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => RESET, Q 
                           => OUT2_24_port, QN => n_2072);
   OUT2_reg_23_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => RESET, Q 
                           => OUT2_23_port, QN => n_2073);
   OUT2_reg_22_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => RESET, Q 
                           => OUT2_22_port, QN => n_2074);
   OUT2_reg_21_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => RESET, Q 
                           => OUT2_21_port, QN => n_2075);
   OUT2_reg_20_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => RESET, Q 
                           => OUT2_20_port, QN => n_2076);
   OUT2_reg_19_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => RESET, Q 
                           => OUT2_19_port, QN => n_2077);
   OUT2_reg_18_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => RESET, Q 
                           => OUT2_18_port, QN => n_2078);
   OUT2_reg_17_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => RESET, Q 
                           => OUT2_17_port, QN => n_2079);
   OUT2_reg_16_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => RESET, Q 
                           => OUT2_16_port, QN => n_2080);
   OUT2_reg_15_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => RESET, Q 
                           => OUT2_15_port, QN => n_2081);
   OUT2_reg_14_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => RESET, Q 
                           => OUT2_14_port, QN => n_2082);
   OUT2_reg_13_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => RESET, Q 
                           => OUT2_13_port, QN => n_2083);
   OUT2_reg_12_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => RESET, Q 
                           => OUT2_12_port, QN => n_2084);
   OUT2_reg_11_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => RESET, Q 
                           => OUT2_11_port, QN => n_2085);
   OUT2_reg_10_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => RESET, Q 
                           => OUT2_10_port, QN => n_2086);
   OUT2_reg_9_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => RESET, Q =>
                           OUT2_9_port, QN => n_2087);
   OUT2_reg_8_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => RESET, Q =>
                           OUT2_8_port, QN => n_2088);
   OUT2_reg_7_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => RESET, Q =>
                           OUT2_7_port, QN => n_2089);
   OUT2_reg_6_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => RESET, Q =>
                           OUT2_6_port, QN => n_2090);
   OUT2_reg_5_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => RESET, Q =>
                           OUT2_5_port, QN => n_2091);
   OUT2_reg_4_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => RESET, Q =>
                           OUT2_4_port, QN => n_2092);
   OUT2_reg_3_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => RESET, Q =>
                           OUT2_3_port, QN => n_2093);
   OUT2_reg_2_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => RESET, Q =>
                           OUT2_2_port, QN => n_2094);
   OUT2_reg_1_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => RESET, Q =>
                           OUT2_1_port, QN => n_2095);
   OUT2_reg_0_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => RESET, Q =>
                           OUT2_0_port, QN => n_2096);
   U2 : NOR2_X1 port map( A1 => n7116, A2 => n7117, ZN => n5332);
   U3 : OR3_X1 port map( A1 => n5293, A2 => n5290, A3 => n5292, ZN => n7116);
   U4 : OR3_X1 port map( A1 => n5289, A2 => n6603, A3 => n5288, ZN => n7117);
   U5 : NOR2_X1 port map( A1 => n7118, A2 => n7119, ZN => n4430);
   U6 : OR3_X1 port map( A1 => n4391, A2 => n4388, A3 => n4390, ZN => n7118);
   U7 : OR3_X1 port map( A1 => n4387, A2 => n6603, A3 => n4386, ZN => n7119);
   U8 : AND2_X1 port map( A1 => n2307, A2 => ADD_WR(1), ZN => n1658);
   U9 : AND2_X1 port map( A1 => n2341, A2 => ADD_WR(1), ZN => n1624);
   U10 : AND2_X1 port map( A1 => n5353, A2 => ADD_WR(1), ZN => n1590);
   U11 : AND2_X1 port map( A1 => n2419, A2 => ADD_WR(1), ZN => n1555);
   U12 : NAND4_X1 port map( A1 => n5300, A2 => n5301, A3 => n5302, A4 => n5303,
                           ZN => n5276);
   U13 : NAND4_X1 port map( A1 => n5258, A2 => n5259, A3 => n5260, A4 => n5261,
                           ZN => n5250);
   U14 : NAND4_X1 port map( A1 => n5232, A2 => n5233, A3 => n5234, A4 => n5235,
                           ZN => n5224);
   U15 : NAND4_X1 port map( A1 => n5206, A2 => n5207, A3 => n5208, A4 => n5209,
                           ZN => n5198);
   U16 : NAND4_X1 port map( A1 => n5180, A2 => n5181, A3 => n5182, A4 => n5183,
                           ZN => n5172);
   U17 : NAND4_X1 port map( A1 => n5154, A2 => n5155, A3 => n5156, A4 => n5157,
                           ZN => n5146);
   U18 : NAND4_X1 port map( A1 => n5128, A2 => n5129, A3 => n5130, A4 => n5131,
                           ZN => n5120);
   U19 : NAND4_X1 port map( A1 => n5102, A2 => n5103, A3 => n5104, A4 => n5105,
                           ZN => n5094);
   U22 : NAND4_X1 port map( A1 => n5076, A2 => n5077, A3 => n5078, A4 => n5079,
                           ZN => n5068);
   U23 : NAND4_X1 port map( A1 => n5050, A2 => n5051, A3 => n5052, A4 => n5053,
                           ZN => n5042);
   U26 : NAND4_X1 port map( A1 => n5024, A2 => n5025, A3 => n5026, A4 => n5027,
                           ZN => n5016);
   U27 : NAND4_X1 port map( A1 => n4998, A2 => n4999, A3 => n5000, A4 => n5001,
                           ZN => n4990);
   U28 : NAND4_X1 port map( A1 => n4972, A2 => n4973, A3 => n4974, A4 => n4975,
                           ZN => n4964);
   U29 : NAND4_X1 port map( A1 => n4946, A2 => n4947, A3 => n4948, A4 => n4949,
                           ZN => n4938);
   U30 : NAND4_X1 port map( A1 => n4920, A2 => n4921, A3 => n4922, A4 => n4923,
                           ZN => n4912);
   U31 : NAND4_X1 port map( A1 => n4894, A2 => n4895, A3 => n4896, A4 => n4897,
                           ZN => n4886);
   U32 : NAND4_X1 port map( A1 => n4868, A2 => n4869, A3 => n4870, A4 => n4871,
                           ZN => n4860);
   U33 : NAND4_X1 port map( A1 => n4842, A2 => n4843, A3 => n4844, A4 => n4845,
                           ZN => n4834);
   U35 : NAND4_X1 port map( A1 => n4816, A2 => n4817, A3 => n4818, A4 => n4819,
                           ZN => n4808);
   U36 : NAND4_X1 port map( A1 => n4790, A2 => n4791, A3 => n4792, A4 => n4793,
                           ZN => n4782);
   U38 : NAND4_X1 port map( A1 => n4764, A2 => n4765, A3 => n4766, A4 => n4767,
                           ZN => n4756);
   U39 : NAND4_X1 port map( A1 => n4738, A2 => n4739, A3 => n4740, A4 => n4741,
                           ZN => n4730);
   U40 : NAND4_X1 port map( A1 => n4712, A2 => n4713, A3 => n4714, A4 => n4715,
                           ZN => n4704);
   U41 : NAND4_X1 port map( A1 => n4686, A2 => n4687, A3 => n4688, A4 => n4689,
                           ZN => n4678);
   U42 : NAND4_X1 port map( A1 => n4660, A2 => n4661, A3 => n4662, A4 => n4663,
                           ZN => n4652);
   U43 : NAND4_X1 port map( A1 => n4634, A2 => n4635, A3 => n4636, A4 => n4637,
                           ZN => n4626);
   U44 : NAND4_X1 port map( A1 => n4608, A2 => n4609, A3 => n4610, A4 => n4611,
                           ZN => n4600);
   U45 : NAND4_X1 port map( A1 => n4582, A2 => n4583, A3 => n4584, A4 => n4585,
                           ZN => n4574);
   U46 : NAND4_X1 port map( A1 => n4556, A2 => n4557, A3 => n4558, A4 => n4559,
                           ZN => n4548);
   U48 : NAND4_X1 port map( A1 => n4530, A2 => n4531, A3 => n4532, A4 => n4533,
                           ZN => n4522);
   U49 : NAND4_X1 port map( A1 => n4504, A2 => n4505, A3 => n4506, A4 => n4507,
                           ZN => n4496);
   U50 : NAND4_X1 port map( A1 => n4455, A2 => n4456, A3 => n4457, A4 => n4458,
                           ZN => n4438);
   U51 : NAND4_X1 port map( A1 => n4398, A2 => n4399, A3 => n4400, A4 => n4401,
                           ZN => n4374);
   U53 : NAND4_X1 port map( A1 => n4356, A2 => n4357, A3 => n4358, A4 => n4359,
                           ZN => n4348);
   U55 : NAND4_X1 port map( A1 => n4330, A2 => n4331, A3 => n4332, A4 => n4333,
                           ZN => n4322);
   U56 : NAND4_X1 port map( A1 => n4304, A2 => n4305, A3 => n4306, A4 => n4307,
                           ZN => n4296);
   U57 : NAND4_X1 port map( A1 => n4278, A2 => n4279, A3 => n4280, A4 => n4281,
                           ZN => n4270);
   U59 : NAND4_X1 port map( A1 => n4252, A2 => n4253, A3 => n4254, A4 => n4255,
                           ZN => n4244);
   U60 : NAND4_X1 port map( A1 => n4226, A2 => n4227, A3 => n4228, A4 => n4229,
                           ZN => n4218);
   U61 : NAND4_X1 port map( A1 => n4200, A2 => n4201, A3 => n4202, A4 => n4203,
                           ZN => n4192);
   U62 : NAND4_X1 port map( A1 => n3982, A2 => n3983, A3 => n3984, A4 => n3985,
                           ZN => n3974);
   U63 : NAND4_X1 port map( A1 => n3956, A2 => n3957, A3 => n3958, A4 => n3959,
                           ZN => n3948);
   U64 : NAND4_X1 port map( A1 => n3930, A2 => n3931, A3 => n3932, A4 => n3933,
                           ZN => n3922);
   U65 : NAND4_X1 port map( A1 => n3040, A2 => n3041, A3 => n3042, A4 => n3043,
                           ZN => n3032);
   U66 : NAND4_X1 port map( A1 => n3014, A2 => n3015, A3 => n3016, A4 => n3017,
                           ZN => n3006);
   U67 : NAND4_X1 port map( A1 => n2988, A2 => n2989, A3 => n2990, A4 => n2991,
                           ZN => n2980);
   U68 : NAND4_X1 port map( A1 => n2962, A2 => n2963, A3 => n2964, A4 => n2965,
                           ZN => n2954);
   U69 : NAND4_X1 port map( A1 => n2936, A2 => n2937, A3 => n2938, A4 => n2939,
                           ZN => n2928);
   U70 : NAND4_X1 port map( A1 => n2910, A2 => n2911, A3 => n2912, A4 => n2913,
                           ZN => n2902);
   U71 : NAND4_X1 port map( A1 => n2884, A2 => n2885, A3 => n2886, A4 => n2887,
                           ZN => n2876);
   U73 : NAND4_X1 port map( A1 => n2858, A2 => n2859, A3 => n2860, A4 => n2861,
                           ZN => n2850);
   U74 : NAND4_X1 port map( A1 => n2832, A2 => n2833, A3 => n2834, A4 => n2835,
                           ZN => n2800);
   U75 : NAND4_X1 port map( A1 => n2782, A2 => n2783, A3 => n2784, A4 => n2785,
                           ZN => n2774);
   U76 : NAND4_X1 port map( A1 => n2756, A2 => n2757, A3 => n2758, A4 => n2759,
                           ZN => n2748);
   U77 : NAND4_X1 port map( A1 => n2730, A2 => n2731, A3 => n2732, A4 => n2733,
                           ZN => n2722);
   U78 : NAND4_X1 port map( A1 => n2704, A2 => n2705, A3 => n2706, A4 => n2707,
                           ZN => n2696);
   U80 : NAND4_X1 port map( A1 => n2678, A2 => n2679, A3 => n2680, A4 => n2681,
                           ZN => n2670);
   U81 : NAND4_X1 port map( A1 => n2652, A2 => n2653, A3 => n2654, A4 => n2655,
                           ZN => n2644);
   U82 : NAND4_X1 port map( A1 => n2626, A2 => n2627, A3 => n2628, A4 => n2629,
                           ZN => n2618);
   U85 : NAND4_X1 port map( A1 => n2600, A2 => n2601, A3 => n2602, A4 => n2603,
                           ZN => n2592);
   U86 : NAND4_X1 port map( A1 => n2574, A2 => n2575, A3 => n2576, A4 => n2577,
                           ZN => n2566);
   U87 : NAND4_X1 port map( A1 => n2548, A2 => n2549, A3 => n2550, A4 => n2551,
                           ZN => n2540);
   U88 : NAND4_X1 port map( A1 => n2522, A2 => n2523, A3 => n2524, A4 => n2525,
                           ZN => n2514);
   U89 : NAND4_X1 port map( A1 => n2473, A2 => n2474, A3 => n2475, A4 => n2476,
                           ZN => n2456);

end SYN_INTEGER;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N5_0 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 downto 
         0);  data_out : out std_logic_vector (4 downto 0));

end gen_reg_N5_0;

architecture SYN_behav of gen_reg_N5_0 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
      n26 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n22, B2 => n16, A => n21, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n16, A2 => data_in(0), ZN => n21);
   U4 : OAI21_X1 port map( B1 => n23, B2 => n16, A => n20, ZN => n4);
   U5 : NAND2_X1 port map( A1 => data_in(1), A2 => n16, ZN => n20);
   U6 : OAI21_X1 port map( B1 => n24, B2 => n16, A => n19, ZN => n3);
   U7 : NAND2_X1 port map( A1 => data_in(2), A2 => n16, ZN => n19);
   U8 : OAI21_X1 port map( B1 => n25, B2 => n16, A => n18, ZN => n2);
   U9 : NAND2_X1 port map( A1 => data_in(3), A2 => n16, ZN => n18);
   U10 : OAI21_X1 port map( B1 => n26, B2 => n16, A => n17, ZN => n1);
   U11 : NAND2_X1 port map( A1 => data_in(4), A2 => n16, ZN => n17);
   U12 : CLKBUF_X1 port map( A => ld, Z => n16);
   data_out_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           data_out(4), QN => n26);
   data_out_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           data_out(3), QN => n25);
   data_out_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           data_out(2), QN => n24);
   data_out_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           data_out(1), QN => n23);
   data_out_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           data_out(0), QN => n22);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_8 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_8;

architecture SYN_behav of gen_reg_N32_8 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n97, n98, n110, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n174, B2 => n110, A => n147, ZN => n9);
   U3 : NAND2_X1 port map( A1 => ld, A2 => data_in(26), ZN => n147);
   U4 : OAI21_X1 port map( B1 => n175, B2 => n110, A => n146, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(27), A2 => n97, ZN => n146);
   U6 : OAI21_X1 port map( B1 => n176, B2 => n110, A => n145, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(28), A2 => n97, ZN => n145);
   U8 : OAI21_X1 port map( B1 => n177, B2 => n98, A => n144, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(29), A2 => n110, ZN => n144);
   U10 : OAI21_X1 port map( B1 => n178, B2 => n110, A => n143, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(30), A2 => n97, ZN => n143);
   U12 : OAI21_X1 port map( B1 => n179, B2 => n110, A => n142, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(31), A2 => n97, ZN => n142);
   U14 : OAI21_X1 port map( B1 => n148, B2 => n110, A => n141, ZN => n35);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => n98, ZN => n141);
   U16 : OAI21_X1 port map( B1 => n149, B2 => n110, A => n140, ZN => n34);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n98, ZN => n140);
   U18 : OAI21_X1 port map( B1 => n150, B2 => n110, A => n139, ZN => n33);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n97, ZN => n139);
   U20 : OAI21_X1 port map( B1 => n151, B2 => n98, A => n138, ZN => n32);
   U21 : NAND2_X1 port map( A1 => data_in(3), A2 => n110, ZN => n138);
   U22 : OAI21_X1 port map( B1 => n152, B2 => n97, A => n137, ZN => n31);
   U23 : NAND2_X1 port map( A1 => data_in(4), A2 => n98, ZN => n137);
   U24 : OAI21_X1 port map( B1 => n153, B2 => n110, A => n136, ZN => n30);
   U25 : NAND2_X1 port map( A1 => data_in(5), A2 => n97, ZN => n136);
   U26 : OAI21_X1 port map( B1 => n154, B2 => n110, A => n135, ZN => n29);
   U27 : NAND2_X1 port map( A1 => data_in(6), A2 => n98, ZN => n135);
   U28 : OAI21_X1 port map( B1 => n155, B2 => n98, A => n134, ZN => n28);
   U29 : NAND2_X1 port map( A1 => data_in(7), A2 => n97, ZN => n134);
   U30 : OAI21_X1 port map( B1 => n156, B2 => n97, A => n133, ZN => n27);
   U31 : NAND2_X1 port map( A1 => data_in(8), A2 => n98, ZN => n133);
   U32 : OAI21_X1 port map( B1 => n157, B2 => n97, A => n132, ZN => n26);
   U33 : NAND2_X1 port map( A1 => data_in(9), A2 => n98, ZN => n132);
   U34 : OAI21_X1 port map( B1 => n158, B2 => n98, A => n131, ZN => n25);
   U35 : NAND2_X1 port map( A1 => data_in(10), A2 => n98, ZN => n131);
   U36 : OAI21_X1 port map( B1 => n159, B2 => n110, A => n130, ZN => n24);
   U37 : NAND2_X1 port map( A1 => data_in(11), A2 => n110, ZN => n130);
   U38 : OAI21_X1 port map( B1 => n160, B2 => n98, A => n129, ZN => n23);
   U39 : NAND2_X1 port map( A1 => data_in(12), A2 => n98, ZN => n129);
   U40 : OAI21_X1 port map( B1 => n161, B2 => n110, A => n128, ZN => n22);
   U41 : NAND2_X1 port map( A1 => data_in(13), A2 => n97, ZN => n128);
   U42 : OAI21_X1 port map( B1 => n162, B2 => n110, A => n127, ZN => n21);
   U43 : NAND2_X1 port map( A1 => data_in(14), A2 => n98, ZN => n127);
   U44 : OAI21_X1 port map( B1 => n163, B2 => n97, A => n126, ZN => n20);
   U45 : NAND2_X1 port map( A1 => data_in(15), A2 => n97, ZN => n126);
   U46 : OAI21_X1 port map( B1 => n164, B2 => n110, A => n125, ZN => n19);
   U47 : NAND2_X1 port map( A1 => data_in(16), A2 => n98, ZN => n125);
   U48 : OAI21_X1 port map( B1 => n165, B2 => n97, A => n124, ZN => n18);
   U49 : NAND2_X1 port map( A1 => data_in(17), A2 => n97, ZN => n124);
   U50 : OAI21_X1 port map( B1 => n166, B2 => n97, A => n123, ZN => n17);
   U51 : NAND2_X1 port map( A1 => data_in(18), A2 => n98, ZN => n123);
   U52 : OAI21_X1 port map( B1 => n167, B2 => n98, A => n122, ZN => n16);
   U53 : NAND2_X1 port map( A1 => data_in(19), A2 => n97, ZN => n122);
   U54 : OAI21_X1 port map( B1 => n168, B2 => n110, A => n121, ZN => n15);
   U55 : NAND2_X1 port map( A1 => data_in(20), A2 => n98, ZN => n121);
   U56 : OAI21_X1 port map( B1 => n169, B2 => n110, A => n120, ZN => n14);
   U57 : NAND2_X1 port map( A1 => data_in(21), A2 => n97, ZN => n120);
   U58 : OAI21_X1 port map( B1 => n170, B2 => ld, A => n119, ZN => n13);
   U59 : NAND2_X1 port map( A1 => data_in(22), A2 => n98, ZN => n119);
   U60 : OAI21_X1 port map( B1 => n171, B2 => ld, A => n118, ZN => n12);
   U61 : NAND2_X1 port map( A1 => data_in(23), A2 => n97, ZN => n118);
   U62 : OAI21_X1 port map( B1 => n172, B2 => n110, A => n117, ZN => n11);
   U63 : NAND2_X1 port map( A1 => data_in(24), A2 => n98, ZN => n117);
   U64 : OAI21_X1 port map( B1 => n173, B2 => n97, A => n116, ZN => n10);
   U65 : NAND2_X1 port map( A1 => data_in(25), A2 => n98, ZN => n116);
   U70 : CLKBUF_X1 port map( A => ld, Z => n97);
   U71 : CLKBUF_X1 port map( A => ld, Z => n98);
   U82 : CLKBUF_X1 port map( A => ld, Z => n110);
   data_out_reg_31_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n179);
   data_out_reg_30_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n178);
   data_out_reg_29_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n177);
   data_out_reg_28_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n176);
   data_out_reg_27_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n175);
   data_out_reg_26_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n174);
   data_out_reg_25_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(25), QN => n173);
   data_out_reg_24_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(24), QN => n172);
   data_out_reg_23_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(23), QN => n171);
   data_out_reg_22_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n170);
   data_out_reg_21_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n169);
   data_out_reg_20_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n168);
   data_out_reg_19_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n167);
   data_out_reg_18_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n166);
   data_out_reg_17_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n165);
   data_out_reg_16_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n164);
   data_out_reg_15_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n163);
   data_out_reg_14_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n162);
   data_out_reg_13_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n161);
   data_out_reg_12_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n160);
   data_out_reg_11_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n159);
   data_out_reg_10_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n158);
   data_out_reg_9_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n157);
   data_out_reg_8_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n156);
   data_out_reg_7_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n155);
   data_out_reg_6_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n154);
   data_out_reg_5_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n153);
   data_out_reg_4_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n152);
   data_out_reg_3_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n151);
   data_out_reg_2_inst : DFFR_X1 port map( D => n33, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n150);
   data_out_reg_1_inst : DFFR_X1 port map( D => n34, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n149);
   data_out_reg_0_inst : DFFR_X1 port map( D => n35, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n148);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity pc_add_N32_OP24 is

   port( data_in : in std_logic_vector (31 downto 0);  data_out : out 
         std_logic_vector (31 downto 0));

end pc_add_N32_OP24;

architecture SYN_behav of pc_add_N32_OP24 is

   component pc_add_N32_OP24_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n4, n5, n6, n_2097 : std_logic;

begin
   
   n4 <= '0';
   n5 <= '1';
   n6 <= '0';
   add_21 : pc_add_N32_OP24_DW01_add_0 port map( A(31) => data_in(31), A(30) =>
                           data_in(30), A(29) => data_in(29), A(28) => 
                           data_in(28), A(27) => data_in(27), A(26) => 
                           data_in(26), A(25) => data_in(25), A(24) => 
                           data_in(24), A(23) => data_in(23), A(22) => 
                           data_in(22), A(21) => data_in(21), A(20) => 
                           data_in(20), A(19) => data_in(19), A(18) => 
                           data_in(18), A(17) => data_in(17), A(16) => 
                           data_in(16), A(15) => data_in(15), A(14) => 
                           data_in(14), A(13) => data_in(13), A(12) => 
                           data_in(12), A(11) => data_in(11), A(10) => 
                           data_in(10), A(9) => data_in(9), A(8) => data_in(8),
                           A(7) => data_in(7), A(6) => data_in(6), A(5) => 
                           data_in(5), A(4) => data_in(4), A(3) => data_in(3), 
                           A(2) => data_in(2), A(1) => data_in(1), A(0) => 
                           data_in(0), B(31) => n4, B(30) => n4, B(29) => n4, 
                           B(28) => n4, B(27) => n4, B(26) => n4, B(25) => n4, 
                           B(24) => n4, B(23) => n4, B(22) => n4, B(21) => n4, 
                           B(20) => n4, B(19) => n4, B(18) => n4, B(17) => n4, 
                           B(16) => n4, B(15) => n4, B(14) => n4, B(13) => n4, 
                           B(12) => n4, B(11) => n4, B(10) => n4, B(9) => n4, 
                           B(8) => n4, B(7) => n4, B(6) => n4, B(5) => n4, B(4)
                           => n4, B(3) => n4, B(2) => n5, B(1) => n4, B(0) => 
                           n4, CI => n6, SUM(31) => data_out(31), SUM(30) => 
                           data_out(30), SUM(29) => data_out(29), SUM(28) => 
                           data_out(28), SUM(27) => data_out(27), SUM(26) => 
                           data_out(26), SUM(25) => data_out(25), SUM(24) => 
                           data_out(24), SUM(23) => data_out(23), SUM(22) => 
                           data_out(22), SUM(21) => data_out(21), SUM(20) => 
                           data_out(20), SUM(19) => data_out(19), SUM(18) => 
                           data_out(18), SUM(17) => data_out(17), SUM(16) => 
                           data_out(16), SUM(15) => data_out(15), SUM(14) => 
                           data_out(14), SUM(13) => data_out(13), SUM(12) => 
                           data_out(12), SUM(11) => data_out(11), SUM(10) => 
                           data_out(10), SUM(9) => data_out(9), SUM(8) => 
                           data_out(8), SUM(7) => data_out(7), SUM(6) => 
                           data_out(6), SUM(5) => data_out(5), SUM(4) => 
                           data_out(4), SUM(3) => data_out(3), SUM(2) => 
                           data_out(2), SUM(1) => data_out(1), SUM(0) => 
                           data_out(0), CO => n_2097);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity gen_reg_N32_0 is

   port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 downto
         0);  data_out : out std_logic_vector (31 downto 0));

end gen_reg_N32_0;

architecture SYN_behav of gen_reg_N32_0 is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n99, n101, n106, n107, n108, n109, n110, n111, n112, n113, n114
      , n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n161, B2 => ld, A => n137, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n99, A2 => data_in(23), ZN => n137);
   U4 : OAI21_X1 port map( B1 => n162, B2 => ld, A => n136, ZN => n8);
   U5 : NAND2_X1 port map( A1 => data_in(24), A2 => n99, ZN => n136);
   U6 : OAI21_X1 port map( B1 => n163, B2 => n101, A => n135, ZN => n7);
   U7 : NAND2_X1 port map( A1 => data_in(25), A2 => n99, ZN => n135);
   U8 : OAI21_X1 port map( B1 => n164, B2 => n101, A => n134, ZN => n6);
   U9 : NAND2_X1 port map( A1 => data_in(26), A2 => n99, ZN => n134);
   U10 : OAI21_X1 port map( B1 => n165, B2 => n101, A => n133, ZN => n5);
   U11 : NAND2_X1 port map( A1 => data_in(27), A2 => n99, ZN => n133);
   U12 : OAI21_X1 port map( B1 => n166, B2 => ld, A => n132, ZN => n4);
   U13 : NAND2_X1 port map( A1 => data_in(28), A2 => n99, ZN => n132);
   U14 : OAI21_X1 port map( B1 => n138, B2 => n101, A => n131, ZN => n32);
   U15 : NAND2_X1 port map( A1 => data_in(0), A2 => n99, ZN => n131);
   U16 : OAI21_X1 port map( B1 => n139, B2 => n101, A => n130, ZN => n31);
   U17 : NAND2_X1 port map( A1 => data_in(1), A2 => n101, ZN => n130);
   U18 : OAI21_X1 port map( B1 => n140, B2 => ld, A => n129, ZN => n30);
   U19 : NAND2_X1 port map( A1 => data_in(2), A2 => n99, ZN => n129);
   U20 : OAI21_X1 port map( B1 => n167, B2 => n101, A => n128, ZN => n3);
   U21 : NAND2_X1 port map( A1 => data_in(29), A2 => n99, ZN => n128);
   U22 : OAI21_X1 port map( B1 => n141, B2 => n99, A => n127, ZN => n29);
   U23 : NAND2_X1 port map( A1 => data_in(3), A2 => n99, ZN => n127);
   U24 : OAI21_X1 port map( B1 => n142, B2 => n99, A => n126, ZN => n28);
   U25 : NAND2_X1 port map( A1 => data_in(4), A2 => n99, ZN => n126);
   U26 : OAI21_X1 port map( B1 => n143, B2 => ld, A => n125, ZN => n27);
   U27 : NAND2_X1 port map( A1 => data_in(5), A2 => n101, ZN => n125);
   U28 : OAI21_X1 port map( B1 => n144, B2 => n99, A => n124, ZN => n26);
   U29 : NAND2_X1 port map( A1 => data_in(6), A2 => ld, ZN => n124);
   U30 : OAI21_X1 port map( B1 => n145, B2 => n99, A => n123, ZN => n25);
   U31 : NAND2_X1 port map( A1 => data_in(7), A2 => ld, ZN => n123);
   U32 : OAI21_X1 port map( B1 => n146, B2 => ld, A => n122, ZN => n24);
   U33 : NAND2_X1 port map( A1 => data_in(8), A2 => n99, ZN => n122);
   U34 : OAI21_X1 port map( B1 => n147, B2 => ld, A => n121, ZN => n23);
   U35 : NAND2_X1 port map( A1 => data_in(9), A2 => n101, ZN => n121);
   U36 : OAI21_X1 port map( B1 => n148, B2 => ld, A => n120, ZN => n22);
   U37 : NAND2_X1 port map( A1 => data_in(10), A2 => n99, ZN => n120);
   U38 : OAI21_X1 port map( B1 => n149, B2 => ld, A => n119, ZN => n21);
   U39 : NAND2_X1 port map( A1 => data_in(11), A2 => n101, ZN => n119);
   U40 : OAI21_X1 port map( B1 => n150, B2 => ld, A => n118, ZN => n20);
   U41 : NAND2_X1 port map( A1 => data_in(12), A2 => ld, ZN => n118);
   U42 : OAI21_X1 port map( B1 => n168, B2 => ld, A => n117, ZN => n2);
   U43 : NAND2_X1 port map( A1 => data_in(30), A2 => ld, ZN => n117);
   U44 : OAI21_X1 port map( B1 => n151, B2 => n101, A => n116, ZN => n19);
   U45 : NAND2_X1 port map( A1 => data_in(13), A2 => ld, ZN => n116);
   U46 : OAI21_X1 port map( B1 => n152, B2 => ld, A => n115, ZN => n18);
   U47 : NAND2_X1 port map( A1 => data_in(14), A2 => ld, ZN => n115);
   U48 : OAI21_X1 port map( B1 => n153, B2 => n101, A => n114, ZN => n17);
   U49 : NAND2_X1 port map( A1 => data_in(15), A2 => ld, ZN => n114);
   U50 : OAI21_X1 port map( B1 => n154, B2 => n101, A => n113, ZN => n16);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => ld, ZN => n113);
   U52 : OAI21_X1 port map( B1 => n155, B2 => n101, A => n112, ZN => n15);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => ld, ZN => n112);
   U54 : OAI21_X1 port map( B1 => n156, B2 => n101, A => n111, ZN => n14);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => ld, ZN => n111);
   U56 : OAI21_X1 port map( B1 => n157, B2 => n101, A => n110, ZN => n13);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => ld, ZN => n110);
   U58 : OAI21_X1 port map( B1 => n158, B2 => n101, A => n109, ZN => n12);
   U59 : NAND2_X1 port map( A1 => data_in(20), A2 => n99, ZN => n109);
   U60 : OAI21_X1 port map( B1 => n159, B2 => n101, A => n108, ZN => n11);
   U61 : NAND2_X1 port map( A1 => data_in(21), A2 => n99, ZN => n108);
   U62 : OAI21_X1 port map( B1 => n160, B2 => n101, A => n107, ZN => n10);
   U63 : NAND2_X1 port map( A1 => data_in(22), A2 => ld, ZN => n107);
   U64 : OAI21_X1 port map( B1 => n169, B2 => n101, A => n106, ZN => n1);
   U65 : NAND2_X1 port map( A1 => data_in(31), A2 => n99, ZN => n106);
   U71 : CLKBUF_X1 port map( A => ld, Z => n99);
   U72 : CLKBUF_X1 port map( A => ld, Z => n101);
   data_out_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q =>
                           data_out(31), QN => n169);
   data_out_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q =>
                           data_out(30), QN => n168);
   data_out_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q =>
                           data_out(29), QN => n167);
   data_out_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q =>
                           data_out(28), QN => n166);
   data_out_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q =>
                           data_out(27), QN => n165);
   data_out_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q =>
                           data_out(26), QN => n164);
   data_out_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q =>
                           data_out(25), QN => n163);
   data_out_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q =>
                           data_out(24), QN => n162);
   data_out_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q =>
                           data_out(23), QN => n161);
   data_out_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q 
                           => data_out(22), QN => n160);
   data_out_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q 
                           => data_out(21), QN => n159);
   data_out_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q 
                           => data_out(20), QN => n158);
   data_out_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q 
                           => data_out(19), QN => n157);
   data_out_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q 
                           => data_out(18), QN => n156);
   data_out_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q 
                           => data_out(17), QN => n155);
   data_out_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q 
                           => data_out(16), QN => n154);
   data_out_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q 
                           => data_out(15), QN => n153);
   data_out_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q 
                           => data_out(14), QN => n152);
   data_out_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q 
                           => data_out(13), QN => n151);
   data_out_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q 
                           => data_out(12), QN => n150);
   data_out_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q 
                           => data_out(11), QN => n149);
   data_out_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q 
                           => data_out(10), QN => n148);
   data_out_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q =>
                           data_out(9), QN => n147);
   data_out_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q =>
                           data_out(8), QN => n146);
   data_out_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q =>
                           data_out(7), QN => n145);
   data_out_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q =>
                           data_out(6), QN => n144);
   data_out_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q =>
                           data_out(5), QN => n143);
   data_out_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q =>
                           data_out(4), QN => n142);
   data_out_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q =>
                           data_out(3), QN => n141);
   data_out_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q =>
                           data_out(2), QN => n140);
   data_out_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q =>
                           data_out(1), QN => n139);
   data_out_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q =>
                           data_out(0), QN => n138);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity WB_STAGE_N_BITS_DATA32_RF_ADDR5 is

   port( CLK, RST, WB_LATCH_EN, JAL_MUX_SEL, WB_MUX_SEL : in std_logic;  IR_IN 
         : in std_logic_vector (4 downto 0);  MUX_IN2, MUX_IN1, MUX_IN0 : in 
         std_logic_vector (31 downto 0);  WRT_OUT : out std_logic_vector (31 
         downto 0);  IR_OUT : out std_logic_vector (4 downto 0));

end WB_STAGE_N_BITS_DATA32_RF_ADDR5;

architecture SYN_STRUCTURAL of WB_STAGE_N_BITS_DATA32_RF_ADDR5 is

   component gen_mux41_N32
      port( sel : in std_logic_vector (1 downto 0);  w, x, y, z : in 
            std_logic_vector (31 downto 0);  m : out std_logic_vector (31 
            downto 0));
   end component;
   
   component gen_reg_N5_1
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 
            downto 0);  data_out : out std_logic_vector (4 downto 0));
   end component;
   
   component gen_reg_N32_1
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal MUX_OUT_31_port, MUX_OUT_30_port, MUX_OUT_29_port, MUX_OUT_28_port, 
      MUX_OUT_27_port, MUX_OUT_26_port, MUX_OUT_25_port, MUX_OUT_24_port, 
      MUX_OUT_23_port, MUX_OUT_22_port, MUX_OUT_21_port, MUX_OUT_20_port, 
      MUX_OUT_19_port, MUX_OUT_18_port, MUX_OUT_17_port, MUX_OUT_16_port, 
      MUX_OUT_15_port, MUX_OUT_14_port, MUX_OUT_13_port, MUX_OUT_12_port, 
      MUX_OUT_11_port, MUX_OUT_10_port, MUX_OUT_9_port, MUX_OUT_8_port, 
      MUX_OUT_7_port, MUX_OUT_6_port, MUX_OUT_5_port, MUX_OUT_4_port, 
      MUX_OUT_3_port, MUX_OUT_2_port, MUX_OUT_1_port, MUX_OUT_0_port : 
      std_logic;

begin
   
   WRT : gen_reg_N32_1 port map( clk => CLK, rst => RST, ld => WB_LATCH_EN, 
                           data_in(31) => MUX_OUT_31_port, data_in(30) => 
                           MUX_OUT_30_port, data_in(29) => MUX_OUT_29_port, 
                           data_in(28) => MUX_OUT_28_port, data_in(27) => 
                           MUX_OUT_27_port, data_in(26) => MUX_OUT_26_port, 
                           data_in(25) => MUX_OUT_25_port, data_in(24) => 
                           MUX_OUT_24_port, data_in(23) => MUX_OUT_23_port, 
                           data_in(22) => MUX_OUT_22_port, data_in(21) => 
                           MUX_OUT_21_port, data_in(20) => MUX_OUT_20_port, 
                           data_in(19) => MUX_OUT_19_port, data_in(18) => 
                           MUX_OUT_18_port, data_in(17) => MUX_OUT_17_port, 
                           data_in(16) => MUX_OUT_16_port, data_in(15) => 
                           MUX_OUT_15_port, data_in(14) => MUX_OUT_14_port, 
                           data_in(13) => MUX_OUT_13_port, data_in(12) => 
                           MUX_OUT_12_port, data_in(11) => MUX_OUT_11_port, 
                           data_in(10) => MUX_OUT_10_port, data_in(9) => 
                           MUX_OUT_9_port, data_in(8) => MUX_OUT_8_port, 
                           data_in(7) => MUX_OUT_7_port, data_in(6) => 
                           MUX_OUT_6_port, data_in(5) => MUX_OUT_5_port, 
                           data_in(4) => MUX_OUT_4_port, data_in(3) => 
                           MUX_OUT_3_port, data_in(2) => MUX_OUT_2_port, 
                           data_in(1) => MUX_OUT_1_port, data_in(0) => 
                           MUX_OUT_0_port, data_out(31) => WRT_OUT(31), 
                           data_out(30) => WRT_OUT(30), data_out(29) => 
                           WRT_OUT(29), data_out(28) => WRT_OUT(28), 
                           data_out(27) => WRT_OUT(27), data_out(26) => 
                           WRT_OUT(26), data_out(25) => WRT_OUT(25), 
                           data_out(24) => WRT_OUT(24), data_out(23) => 
                           WRT_OUT(23), data_out(22) => WRT_OUT(22), 
                           data_out(21) => WRT_OUT(21), data_out(20) => 
                           WRT_OUT(20), data_out(19) => WRT_OUT(19), 
                           data_out(18) => WRT_OUT(18), data_out(17) => 
                           WRT_OUT(17), data_out(16) => WRT_OUT(16), 
                           data_out(15) => WRT_OUT(15), data_out(14) => 
                           WRT_OUT(14), data_out(13) => WRT_OUT(13), 
                           data_out(12) => WRT_OUT(12), data_out(11) => 
                           WRT_OUT(11), data_out(10) => WRT_OUT(10), 
                           data_out(9) => WRT_OUT(9), data_out(8) => WRT_OUT(8)
                           , data_out(7) => WRT_OUT(7), data_out(6) => 
                           WRT_OUT(6), data_out(5) => WRT_OUT(5), data_out(4) 
                           => WRT_OUT(4), data_out(3) => WRT_OUT(3), 
                           data_out(2) => WRT_OUT(2), data_out(1) => WRT_OUT(1)
                           , data_out(0) => WRT_OUT(0));
   IR4 : gen_reg_N5_1 port map( clk => CLK, rst => RST, ld => WB_LATCH_EN, 
                           data_in(4) => IR_IN(4), data_in(3) => IR_IN(3), 
                           data_in(2) => IR_IN(2), data_in(1) => IR_IN(1), 
                           data_in(0) => IR_IN(0), data_out(4) => IR_OUT(4), 
                           data_out(3) => IR_OUT(3), data_out(2) => IR_OUT(2), 
                           data_out(1) => IR_OUT(1), data_out(0) => IR_OUT(0));
   MUX : gen_mux41_N32 port map( sel(1) => JAL_MUX_SEL, sel(0) => WB_MUX_SEL, 
                           w(31) => MUX_IN0(31), w(30) => MUX_IN0(30), w(29) =>
                           MUX_IN0(29), w(28) => MUX_IN0(28), w(27) => 
                           MUX_IN0(27), w(26) => MUX_IN0(26), w(25) => 
                           MUX_IN0(25), w(24) => MUX_IN0(24), w(23) => 
                           MUX_IN0(23), w(22) => MUX_IN0(22), w(21) => 
                           MUX_IN0(21), w(20) => MUX_IN0(20), w(19) => 
                           MUX_IN0(19), w(18) => MUX_IN0(18), w(17) => 
                           MUX_IN0(17), w(16) => MUX_IN0(16), w(15) => 
                           MUX_IN0(15), w(14) => MUX_IN0(14), w(13) => 
                           MUX_IN0(13), w(12) => MUX_IN0(12), w(11) => 
                           MUX_IN0(11), w(10) => MUX_IN0(10), w(9) => 
                           MUX_IN0(9), w(8) => MUX_IN0(8), w(7) => MUX_IN0(7), 
                           w(6) => MUX_IN0(6), w(5) => MUX_IN0(5), w(4) => 
                           MUX_IN0(4), w(3) => MUX_IN0(3), w(2) => MUX_IN0(2), 
                           w(1) => MUX_IN0(1), w(0) => MUX_IN0(0), x(31) => 
                           MUX_IN1(31), x(30) => MUX_IN1(30), x(29) => 
                           MUX_IN1(29), x(28) => MUX_IN1(28), x(27) => 
                           MUX_IN1(27), x(26) => MUX_IN1(26), x(25) => 
                           MUX_IN1(25), x(24) => MUX_IN1(24), x(23) => 
                           MUX_IN1(23), x(22) => MUX_IN1(22), x(21) => 
                           MUX_IN1(21), x(20) => MUX_IN1(20), x(19) => 
                           MUX_IN1(19), x(18) => MUX_IN1(18), x(17) => 
                           MUX_IN1(17), x(16) => MUX_IN1(16), x(15) => 
                           MUX_IN1(15), x(14) => MUX_IN1(14), x(13) => 
                           MUX_IN1(13), x(12) => MUX_IN1(12), x(11) => 
                           MUX_IN1(11), x(10) => MUX_IN1(10), x(9) => 
                           MUX_IN1(9), x(8) => MUX_IN1(8), x(7) => MUX_IN1(7), 
                           x(6) => MUX_IN1(6), x(5) => MUX_IN1(5), x(4) => 
                           MUX_IN1(4), x(3) => MUX_IN1(3), x(2) => MUX_IN1(2), 
                           x(1) => MUX_IN1(1), x(0) => MUX_IN1(0), y(31) => 
                           MUX_IN2(31), y(30) => MUX_IN2(30), y(29) => 
                           MUX_IN2(29), y(28) => MUX_IN2(28), y(27) => 
                           MUX_IN2(27), y(26) => MUX_IN2(26), y(25) => 
                           MUX_IN2(25), y(24) => MUX_IN2(24), y(23) => 
                           MUX_IN2(23), y(22) => MUX_IN2(22), y(21) => 
                           MUX_IN2(21), y(20) => MUX_IN2(20), y(19) => 
                           MUX_IN2(19), y(18) => MUX_IN2(18), y(17) => 
                           MUX_IN2(17), y(16) => MUX_IN2(16), y(15) => 
                           MUX_IN2(15), y(14) => MUX_IN2(14), y(13) => 
                           MUX_IN2(13), y(12) => MUX_IN2(12), y(11) => 
                           MUX_IN2(11), y(10) => MUX_IN2(10), y(9) => 
                           MUX_IN2(9), y(8) => MUX_IN2(8), y(7) => MUX_IN2(7), 
                           y(6) => MUX_IN2(6), y(5) => MUX_IN2(5), y(4) => 
                           MUX_IN2(4), y(3) => MUX_IN2(3), y(2) => MUX_IN2(2), 
                           y(1) => MUX_IN2(1), y(0) => MUX_IN2(0), z(31) => 
                           MUX_IN2(31), z(30) => MUX_IN2(30), z(29) => 
                           MUX_IN2(29), z(28) => MUX_IN2(28), z(27) => 
                           MUX_IN2(27), z(26) => MUX_IN2(26), z(25) => 
                           MUX_IN2(25), z(24) => MUX_IN2(24), z(23) => 
                           MUX_IN2(23), z(22) => MUX_IN2(22), z(21) => 
                           MUX_IN2(21), z(20) => MUX_IN2(20), z(19) => 
                           MUX_IN2(19), z(18) => MUX_IN2(18), z(17) => 
                           MUX_IN2(17), z(16) => MUX_IN2(16), z(15) => 
                           MUX_IN2(15), z(14) => MUX_IN2(14), z(13) => 
                           MUX_IN2(13), z(12) => MUX_IN2(12), z(11) => 
                           MUX_IN2(11), z(10) => MUX_IN2(10), z(9) => 
                           MUX_IN2(9), z(8) => MUX_IN2(8), z(7) => MUX_IN2(7), 
                           z(6) => MUX_IN2(6), z(5) => MUX_IN2(5), z(4) => 
                           MUX_IN2(4), z(3) => MUX_IN2(3), z(2) => MUX_IN2(2), 
                           z(1) => MUX_IN2(1), z(0) => MUX_IN2(0), m(31) => 
                           MUX_OUT_31_port, m(30) => MUX_OUT_30_port, m(29) => 
                           MUX_OUT_29_port, m(28) => MUX_OUT_28_port, m(27) => 
                           MUX_OUT_27_port, m(26) => MUX_OUT_26_port, m(25) => 
                           MUX_OUT_25_port, m(24) => MUX_OUT_24_port, m(23) => 
                           MUX_OUT_23_port, m(22) => MUX_OUT_22_port, m(21) => 
                           MUX_OUT_21_port, m(20) => MUX_OUT_20_port, m(19) => 
                           MUX_OUT_19_port, m(18) => MUX_OUT_18_port, m(17) => 
                           MUX_OUT_17_port, m(16) => MUX_OUT_16_port, m(15) => 
                           MUX_OUT_15_port, m(14) => MUX_OUT_14_port, m(13) => 
                           MUX_OUT_13_port, m(12) => MUX_OUT_12_port, m(11) => 
                           MUX_OUT_11_port, m(10) => MUX_OUT_10_port, m(9) => 
                           MUX_OUT_9_port, m(8) => MUX_OUT_8_port, m(7) => 
                           MUX_OUT_7_port, m(6) => MUX_OUT_6_port, m(5) => 
                           MUX_OUT_5_port, m(4) => MUX_OUT_4_port, m(3) => 
                           MUX_OUT_3_port, m(2) => MUX_OUT_2_port, m(1) => 
                           MUX_OUT_1_port, m(0) => MUX_OUT_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity MEM_STAGE_N_BITS_DATA32_RF_ADDR5 is

   port( CLK, RST, MEM_OUTREG_EN, ZERO_PADDING4, MEM_OUT_SEL : in std_logic;  
         BYTE_LEN_IN : in std_logic_vector (1 downto 0);  DRAM_WE : in 
         std_logic;  DRAM_WE_OUT : out std_logic;  BYTE_LEN_OUT : out 
         std_logic_vector (1 downto 0);  BRA_IN : in std_logic;  JUMP_MUX_IN_0,
         ALU_OUTPUT_IN, MEM_DATA_IN, MEM_DATA_OUT_INT, NPC_IN : in 
         std_logic_vector (31 downto 0);  IR_IN : in std_logic_vector (4 downto
         0);  IR_OUT : out std_logic_vector (4 downto 0);  NPC_OUT, 
         MEM_ADDR_OUT, MEM_DATA_IN_PRIME, ALU_OUTPUT_OUT, MEM_DATA_OUT, 
         ADDR_MUX_OUT : out std_logic_vector (31 downto 0));

end MEM_STAGE_N_BITS_DATA32_RF_ADDR5;

architecture SYN_STRUCTURAL of MEM_STAGE_N_BITS_DATA32_RF_ADDR5 is

   component sign_ext_alt_N_IN016_N_IN18_N_OUT32
      port( ctrl_in, zero_padding : in std_logic;  data_in : in 
            std_logic_vector (15 downto 0);  data_ext : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component gen_reg_N5_2
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 
            downto 0);  data_out : out std_logic_vector (4 downto 0));
   end component;
   
   component gen_reg_N32_2
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N32_3
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N1_1
      port( clk, rst, ld, data_in : in std_logic;  data_out : out std_logic);
   end component;
   
   component gen_mux21_N32_1
      port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m :
            out std_logic_vector (31 downto 0));
   end component;
   
   component gen_mux21_N32_2
      port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal ALU_OUTPUT_OUT_31_port, ALU_OUTPUT_OUT_30_port, 
      ALU_OUTPUT_OUT_29_port, ALU_OUTPUT_OUT_28_port, ALU_OUTPUT_OUT_27_port, 
      ALU_OUTPUT_OUT_26_port, ALU_OUTPUT_OUT_25_port, ALU_OUTPUT_OUT_24_port, 
      ALU_OUTPUT_OUT_23_port, ALU_OUTPUT_OUT_22_port, ALU_OUTPUT_OUT_21_port, 
      ALU_OUTPUT_OUT_20_port, ALU_OUTPUT_OUT_19_port, ALU_OUTPUT_OUT_18_port, 
      ALU_OUTPUT_OUT_17_port, ALU_OUTPUT_OUT_16_port, ALU_OUTPUT_OUT_15_port, 
      ALU_OUTPUT_OUT_14_port, ALU_OUTPUT_OUT_13_port, ALU_OUTPUT_OUT_12_port, 
      ALU_OUTPUT_OUT_11_port, ALU_OUTPUT_OUT_10_port, ALU_OUTPUT_OUT_9_port, 
      ALU_OUTPUT_OUT_8_port, ALU_OUTPUT_OUT_7_port, ALU_OUTPUT_OUT_6_port, 
      ALU_OUTPUT_OUT_5_port, ALU_OUTPUT_OUT_4_port, ALU_OUTPUT_OUT_3_port, 
      ALU_OUTPUT_OUT_2_port, ALU_OUTPUT_OUT_1_port, ALU_OUTPUT_OUT_0_port, 
      BRA_OUT_AUX_0_port, SIGN_EXT_OUT_31_port, SIGN_EXT_OUT_30_port, 
      SIGN_EXT_OUT_29_port, SIGN_EXT_OUT_28_port, SIGN_EXT_OUT_27_port, 
      SIGN_EXT_OUT_26_port, SIGN_EXT_OUT_25_port, SIGN_EXT_OUT_24_port, 
      SIGN_EXT_OUT_23_port, SIGN_EXT_OUT_22_port, SIGN_EXT_OUT_21_port, 
      SIGN_EXT_OUT_20_port, SIGN_EXT_OUT_19_port, SIGN_EXT_OUT_18_port, 
      SIGN_EXT_OUT_17_port, SIGN_EXT_OUT_16_port, SIGN_EXT_OUT_15_port, 
      SIGN_EXT_OUT_14_port, SIGN_EXT_OUT_13_port, SIGN_EXT_OUT_12_port, 
      SIGN_EXT_OUT_11_port, SIGN_EXT_OUT_10_port, SIGN_EXT_OUT_9_port, 
      SIGN_EXT_OUT_8_port, SIGN_EXT_OUT_7_port, SIGN_EXT_OUT_6_port, 
      SIGN_EXT_OUT_5_port, SIGN_EXT_OUT_4_port, SIGN_EXT_OUT_3_port, 
      SIGN_EXT_OUT_2_port, SIGN_EXT_OUT_1_port, SIGN_EXT_OUT_0_port : std_logic
      ;

begin
   DRAM_WE_OUT <= DRAM_WE;
   BYTE_LEN_OUT <= ( BYTE_LEN_IN(1), BYTE_LEN_IN(0) );
   MEM_ADDR_OUT <= ( ALU_OUTPUT_IN(31), ALU_OUTPUT_IN(30), ALU_OUTPUT_IN(29), 
      ALU_OUTPUT_IN(28), ALU_OUTPUT_IN(27), ALU_OUTPUT_IN(26), 
      ALU_OUTPUT_IN(25), ALU_OUTPUT_IN(24), ALU_OUTPUT_IN(23), 
      ALU_OUTPUT_IN(22), ALU_OUTPUT_IN(21), ALU_OUTPUT_IN(20), 
      ALU_OUTPUT_IN(19), ALU_OUTPUT_IN(18), ALU_OUTPUT_IN(17), 
      ALU_OUTPUT_IN(16), ALU_OUTPUT_IN(15), ALU_OUTPUT_IN(14), 
      ALU_OUTPUT_IN(13), ALU_OUTPUT_IN(12), ALU_OUTPUT_IN(11), 
      ALU_OUTPUT_IN(10), ALU_OUTPUT_IN(9), ALU_OUTPUT_IN(8), ALU_OUTPUT_IN(7), 
      ALU_OUTPUT_IN(6), ALU_OUTPUT_IN(5), ALU_OUTPUT_IN(4), ALU_OUTPUT_IN(3), 
      ALU_OUTPUT_IN(2), ALU_OUTPUT_IN(1), ALU_OUTPUT_IN(0) );
   MEM_DATA_IN_PRIME <= ( MEM_DATA_IN(31), MEM_DATA_IN(30), MEM_DATA_IN(29), 
      MEM_DATA_IN(28), MEM_DATA_IN(27), MEM_DATA_IN(26), MEM_DATA_IN(25), 
      MEM_DATA_IN(24), MEM_DATA_IN(23), MEM_DATA_IN(22), MEM_DATA_IN(21), 
      MEM_DATA_IN(20), MEM_DATA_IN(19), MEM_DATA_IN(18), MEM_DATA_IN(17), 
      MEM_DATA_IN(16), MEM_DATA_IN(15), MEM_DATA_IN(14), MEM_DATA_IN(13), 
      MEM_DATA_IN(12), MEM_DATA_IN(11), MEM_DATA_IN(10), MEM_DATA_IN(9), 
      MEM_DATA_IN(8), MEM_DATA_IN(7), MEM_DATA_IN(6), MEM_DATA_IN(5), 
      MEM_DATA_IN(4), MEM_DATA_IN(3), MEM_DATA_IN(2), MEM_DATA_IN(1), 
      MEM_DATA_IN(0) );
   ALU_OUTPUT_OUT <= ( ALU_OUTPUT_OUT_31_port, ALU_OUTPUT_OUT_30_port, 
      ALU_OUTPUT_OUT_29_port, ALU_OUTPUT_OUT_28_port, ALU_OUTPUT_OUT_27_port, 
      ALU_OUTPUT_OUT_26_port, ALU_OUTPUT_OUT_25_port, ALU_OUTPUT_OUT_24_port, 
      ALU_OUTPUT_OUT_23_port, ALU_OUTPUT_OUT_22_port, ALU_OUTPUT_OUT_21_port, 
      ALU_OUTPUT_OUT_20_port, ALU_OUTPUT_OUT_19_port, ALU_OUTPUT_OUT_18_port, 
      ALU_OUTPUT_OUT_17_port, ALU_OUTPUT_OUT_16_port, ALU_OUTPUT_OUT_15_port, 
      ALU_OUTPUT_OUT_14_port, ALU_OUTPUT_OUT_13_port, ALU_OUTPUT_OUT_12_port, 
      ALU_OUTPUT_OUT_11_port, ALU_OUTPUT_OUT_10_port, ALU_OUTPUT_OUT_9_port, 
      ALU_OUTPUT_OUT_8_port, ALU_OUTPUT_OUT_7_port, ALU_OUTPUT_OUT_6_port, 
      ALU_OUTPUT_OUT_5_port, ALU_OUTPUT_OUT_4_port, ALU_OUTPUT_OUT_3_port, 
      ALU_OUTPUT_OUT_2_port, ALU_OUTPUT_OUT_1_port, ALU_OUTPUT_OUT_0_port );
   
   ADDR_MUX : gen_mux21_N32_2 port map( sel => BRA_OUT_AUX_0_port, x(31) => 
                           JUMP_MUX_IN_0(31), x(30) => JUMP_MUX_IN_0(30), x(29)
                           => JUMP_MUX_IN_0(29), x(28) => JUMP_MUX_IN_0(28), 
                           x(27) => JUMP_MUX_IN_0(27), x(26) => 
                           JUMP_MUX_IN_0(26), x(25) => JUMP_MUX_IN_0(25), x(24)
                           => JUMP_MUX_IN_0(24), x(23) => JUMP_MUX_IN_0(23), 
                           x(22) => JUMP_MUX_IN_0(22), x(21) => 
                           JUMP_MUX_IN_0(21), x(20) => JUMP_MUX_IN_0(20), x(19)
                           => JUMP_MUX_IN_0(19), x(18) => JUMP_MUX_IN_0(18), 
                           x(17) => JUMP_MUX_IN_0(17), x(16) => 
                           JUMP_MUX_IN_0(16), x(15) => JUMP_MUX_IN_0(15), x(14)
                           => JUMP_MUX_IN_0(14), x(13) => JUMP_MUX_IN_0(13), 
                           x(12) => JUMP_MUX_IN_0(12), x(11) => 
                           JUMP_MUX_IN_0(11), x(10) => JUMP_MUX_IN_0(10), x(9) 
                           => JUMP_MUX_IN_0(9), x(8) => JUMP_MUX_IN_0(8), x(7) 
                           => JUMP_MUX_IN_0(7), x(6) => JUMP_MUX_IN_0(6), x(5) 
                           => JUMP_MUX_IN_0(5), x(4) => JUMP_MUX_IN_0(4), x(3) 
                           => JUMP_MUX_IN_0(3), x(2) => JUMP_MUX_IN_0(2), x(1) 
                           => JUMP_MUX_IN_0(1), x(0) => JUMP_MUX_IN_0(0), y(31)
                           => ALU_OUTPUT_OUT_31_port, y(30) => 
                           ALU_OUTPUT_OUT_30_port, y(29) => 
                           ALU_OUTPUT_OUT_29_port, y(28) => 
                           ALU_OUTPUT_OUT_28_port, y(27) => 
                           ALU_OUTPUT_OUT_27_port, y(26) => 
                           ALU_OUTPUT_OUT_26_port, y(25) => 
                           ALU_OUTPUT_OUT_25_port, y(24) => 
                           ALU_OUTPUT_OUT_24_port, y(23) => 
                           ALU_OUTPUT_OUT_23_port, y(22) => 
                           ALU_OUTPUT_OUT_22_port, y(21) => 
                           ALU_OUTPUT_OUT_21_port, y(20) => 
                           ALU_OUTPUT_OUT_20_port, y(19) => 
                           ALU_OUTPUT_OUT_19_port, y(18) => 
                           ALU_OUTPUT_OUT_18_port, y(17) => 
                           ALU_OUTPUT_OUT_17_port, y(16) => 
                           ALU_OUTPUT_OUT_16_port, y(15) => 
                           ALU_OUTPUT_OUT_15_port, y(14) => 
                           ALU_OUTPUT_OUT_14_port, y(13) => 
                           ALU_OUTPUT_OUT_13_port, y(12) => 
                           ALU_OUTPUT_OUT_12_port, y(11) => 
                           ALU_OUTPUT_OUT_11_port, y(10) => 
                           ALU_OUTPUT_OUT_10_port, y(9) => 
                           ALU_OUTPUT_OUT_9_port, y(8) => ALU_OUTPUT_OUT_8_port
                           , y(7) => ALU_OUTPUT_OUT_7_port, y(6) => 
                           ALU_OUTPUT_OUT_6_port, y(5) => ALU_OUTPUT_OUT_5_port
                           , y(4) => ALU_OUTPUT_OUT_4_port, y(3) => 
                           ALU_OUTPUT_OUT_3_port, y(2) => ALU_OUTPUT_OUT_2_port
                           , y(1) => ALU_OUTPUT_OUT_1_port, y(0) => 
                           ALU_OUTPUT_OUT_0_port, m(31) => ADDR_MUX_OUT(31), 
                           m(30) => ADDR_MUX_OUT(30), m(29) => ADDR_MUX_OUT(29)
                           , m(28) => ADDR_MUX_OUT(28), m(27) => 
                           ADDR_MUX_OUT(27), m(26) => ADDR_MUX_OUT(26), m(25) 
                           => ADDR_MUX_OUT(25), m(24) => ADDR_MUX_OUT(24), 
                           m(23) => ADDR_MUX_OUT(23), m(22) => ADDR_MUX_OUT(22)
                           , m(21) => ADDR_MUX_OUT(21), m(20) => 
                           ADDR_MUX_OUT(20), m(19) => ADDR_MUX_OUT(19), m(18) 
                           => ADDR_MUX_OUT(18), m(17) => ADDR_MUX_OUT(17), 
                           m(16) => ADDR_MUX_OUT(16), m(15) => ADDR_MUX_OUT(15)
                           , m(14) => ADDR_MUX_OUT(14), m(13) => 
                           ADDR_MUX_OUT(13), m(12) => ADDR_MUX_OUT(12), m(11) 
                           => ADDR_MUX_OUT(11), m(10) => ADDR_MUX_OUT(10), m(9)
                           => ADDR_MUX_OUT(9), m(8) => ADDR_MUX_OUT(8), m(7) =>
                           ADDR_MUX_OUT(7), m(6) => ADDR_MUX_OUT(6), m(5) => 
                           ADDR_MUX_OUT(5), m(4) => ADDR_MUX_OUT(4), m(3) => 
                           ADDR_MUX_OUT(3), m(2) => ADDR_MUX_OUT(2), m(1) => 
                           ADDR_MUX_OUT(1), m(0) => ADDR_MUX_OUT(0));
   DATA_MUX : gen_mux21_N32_1 port map( sel => MEM_OUT_SEL, x(31) => 
                           SIGN_EXT_OUT_31_port, x(30) => SIGN_EXT_OUT_30_port,
                           x(29) => SIGN_EXT_OUT_29_port, x(28) => 
                           SIGN_EXT_OUT_28_port, x(27) => SIGN_EXT_OUT_27_port,
                           x(26) => SIGN_EXT_OUT_26_port, x(25) => 
                           SIGN_EXT_OUT_25_port, x(24) => SIGN_EXT_OUT_24_port,
                           x(23) => SIGN_EXT_OUT_23_port, x(22) => 
                           SIGN_EXT_OUT_22_port, x(21) => SIGN_EXT_OUT_21_port,
                           x(20) => SIGN_EXT_OUT_20_port, x(19) => 
                           SIGN_EXT_OUT_19_port, x(18) => SIGN_EXT_OUT_18_port,
                           x(17) => SIGN_EXT_OUT_17_port, x(16) => 
                           SIGN_EXT_OUT_16_port, x(15) => SIGN_EXT_OUT_15_port,
                           x(14) => SIGN_EXT_OUT_14_port, x(13) => 
                           SIGN_EXT_OUT_13_port, x(12) => SIGN_EXT_OUT_12_port,
                           x(11) => SIGN_EXT_OUT_11_port, x(10) => 
                           SIGN_EXT_OUT_10_port, x(9) => SIGN_EXT_OUT_9_port, 
                           x(8) => SIGN_EXT_OUT_8_port, x(7) => 
                           SIGN_EXT_OUT_7_port, x(6) => SIGN_EXT_OUT_6_port, 
                           x(5) => SIGN_EXT_OUT_5_port, x(4) => 
                           SIGN_EXT_OUT_4_port, x(3) => SIGN_EXT_OUT_3_port, 
                           x(2) => SIGN_EXT_OUT_2_port, x(1) => 
                           SIGN_EXT_OUT_1_port, x(0) => SIGN_EXT_OUT_0_port, 
                           y(31) => MEM_DATA_OUT_INT(31), y(30) => 
                           MEM_DATA_OUT_INT(30), y(29) => MEM_DATA_OUT_INT(29),
                           y(28) => MEM_DATA_OUT_INT(28), y(27) => 
                           MEM_DATA_OUT_INT(27), y(26) => MEM_DATA_OUT_INT(26),
                           y(25) => MEM_DATA_OUT_INT(25), y(24) => 
                           MEM_DATA_OUT_INT(24), y(23) => MEM_DATA_OUT_INT(23),
                           y(22) => MEM_DATA_OUT_INT(22), y(21) => 
                           MEM_DATA_OUT_INT(21), y(20) => MEM_DATA_OUT_INT(20),
                           y(19) => MEM_DATA_OUT_INT(19), y(18) => 
                           MEM_DATA_OUT_INT(18), y(17) => MEM_DATA_OUT_INT(17),
                           y(16) => MEM_DATA_OUT_INT(16), y(15) => 
                           MEM_DATA_OUT_INT(15), y(14) => MEM_DATA_OUT_INT(14),
                           y(13) => MEM_DATA_OUT_INT(13), y(12) => 
                           MEM_DATA_OUT_INT(12), y(11) => MEM_DATA_OUT_INT(11),
                           y(10) => MEM_DATA_OUT_INT(10), y(9) => 
                           MEM_DATA_OUT_INT(9), y(8) => MEM_DATA_OUT_INT(8), 
                           y(7) => MEM_DATA_OUT_INT(7), y(6) => 
                           MEM_DATA_OUT_INT(6), y(5) => MEM_DATA_OUT_INT(5), 
                           y(4) => MEM_DATA_OUT_INT(4), y(3) => 
                           MEM_DATA_OUT_INT(3), y(2) => MEM_DATA_OUT_INT(2), 
                           y(1) => MEM_DATA_OUT_INT(1), y(0) => 
                           MEM_DATA_OUT_INT(0), m(31) => MEM_DATA_OUT(31), 
                           m(30) => MEM_DATA_OUT(30), m(29) => MEM_DATA_OUT(29)
                           , m(28) => MEM_DATA_OUT(28), m(27) => 
                           MEM_DATA_OUT(27), m(26) => MEM_DATA_OUT(26), m(25) 
                           => MEM_DATA_OUT(25), m(24) => MEM_DATA_OUT(24), 
                           m(23) => MEM_DATA_OUT(23), m(22) => MEM_DATA_OUT(22)
                           , m(21) => MEM_DATA_OUT(21), m(20) => 
                           MEM_DATA_OUT(20), m(19) => MEM_DATA_OUT(19), m(18) 
                           => MEM_DATA_OUT(18), m(17) => MEM_DATA_OUT(17), 
                           m(16) => MEM_DATA_OUT(16), m(15) => MEM_DATA_OUT(15)
                           , m(14) => MEM_DATA_OUT(14), m(13) => 
                           MEM_DATA_OUT(13), m(12) => MEM_DATA_OUT(12), m(11) 
                           => MEM_DATA_OUT(11), m(10) => MEM_DATA_OUT(10), m(9)
                           => MEM_DATA_OUT(9), m(8) => MEM_DATA_OUT(8), m(7) =>
                           MEM_DATA_OUT(7), m(6) => MEM_DATA_OUT(6), m(5) => 
                           MEM_DATA_OUT(5), m(4) => MEM_DATA_OUT(4), m(3) => 
                           MEM_DATA_OUT(3), m(2) => MEM_DATA_OUT(2), m(1) => 
                           MEM_DATA_OUT(1), m(0) => MEM_DATA_OUT(0));
   BRA : gen_reg_N1_1 port map( clk => CLK, rst => RST, ld => MEM_OUTREG_EN, 
                           data_in => BRA_IN, data_out => BRA_OUT_AUX_0_port);
   ALU_OUTPUT : gen_reg_N32_3 port map( clk => CLK, rst => RST, ld => 
                           MEM_OUTREG_EN, data_in(31) => ALU_OUTPUT_IN(31), 
                           data_in(30) => ALU_OUTPUT_IN(30), data_in(29) => 
                           ALU_OUTPUT_IN(29), data_in(28) => ALU_OUTPUT_IN(28),
                           data_in(27) => ALU_OUTPUT_IN(27), data_in(26) => 
                           ALU_OUTPUT_IN(26), data_in(25) => ALU_OUTPUT_IN(25),
                           data_in(24) => ALU_OUTPUT_IN(24), data_in(23) => 
                           ALU_OUTPUT_IN(23), data_in(22) => ALU_OUTPUT_IN(22),
                           data_in(21) => ALU_OUTPUT_IN(21), data_in(20) => 
                           ALU_OUTPUT_IN(20), data_in(19) => ALU_OUTPUT_IN(19),
                           data_in(18) => ALU_OUTPUT_IN(18), data_in(17) => 
                           ALU_OUTPUT_IN(17), data_in(16) => ALU_OUTPUT_IN(16),
                           data_in(15) => ALU_OUTPUT_IN(15), data_in(14) => 
                           ALU_OUTPUT_IN(14), data_in(13) => ALU_OUTPUT_IN(13),
                           data_in(12) => ALU_OUTPUT_IN(12), data_in(11) => 
                           ALU_OUTPUT_IN(11), data_in(10) => ALU_OUTPUT_IN(10),
                           data_in(9) => ALU_OUTPUT_IN(9), data_in(8) => 
                           ALU_OUTPUT_IN(8), data_in(7) => ALU_OUTPUT_IN(7), 
                           data_in(6) => ALU_OUTPUT_IN(6), data_in(5) => 
                           ALU_OUTPUT_IN(5), data_in(4) => ALU_OUTPUT_IN(4), 
                           data_in(3) => ALU_OUTPUT_IN(3), data_in(2) => 
                           ALU_OUTPUT_IN(2), data_in(1) => ALU_OUTPUT_IN(1), 
                           data_in(0) => ALU_OUTPUT_IN(0), data_out(31) => 
                           ALU_OUTPUT_OUT_31_port, data_out(30) => 
                           ALU_OUTPUT_OUT_30_port, data_out(29) => 
                           ALU_OUTPUT_OUT_29_port, data_out(28) => 
                           ALU_OUTPUT_OUT_28_port, data_out(27) => 
                           ALU_OUTPUT_OUT_27_port, data_out(26) => 
                           ALU_OUTPUT_OUT_26_port, data_out(25) => 
                           ALU_OUTPUT_OUT_25_port, data_out(24) => 
                           ALU_OUTPUT_OUT_24_port, data_out(23) => 
                           ALU_OUTPUT_OUT_23_port, data_out(22) => 
                           ALU_OUTPUT_OUT_22_port, data_out(21) => 
                           ALU_OUTPUT_OUT_21_port, data_out(20) => 
                           ALU_OUTPUT_OUT_20_port, data_out(19) => 
                           ALU_OUTPUT_OUT_19_port, data_out(18) => 
                           ALU_OUTPUT_OUT_18_port, data_out(17) => 
                           ALU_OUTPUT_OUT_17_port, data_out(16) => 
                           ALU_OUTPUT_OUT_16_port, data_out(15) => 
                           ALU_OUTPUT_OUT_15_port, data_out(14) => 
                           ALU_OUTPUT_OUT_14_port, data_out(13) => 
                           ALU_OUTPUT_OUT_13_port, data_out(12) => 
                           ALU_OUTPUT_OUT_12_port, data_out(11) => 
                           ALU_OUTPUT_OUT_11_port, data_out(10) => 
                           ALU_OUTPUT_OUT_10_port, data_out(9) => 
                           ALU_OUTPUT_OUT_9_port, data_out(8) => 
                           ALU_OUTPUT_OUT_8_port, data_out(7) => 
                           ALU_OUTPUT_OUT_7_port, data_out(6) => 
                           ALU_OUTPUT_OUT_6_port, data_out(5) => 
                           ALU_OUTPUT_OUT_5_port, data_out(4) => 
                           ALU_OUTPUT_OUT_4_port, data_out(3) => 
                           ALU_OUTPUT_OUT_3_port, data_out(2) => 
                           ALU_OUTPUT_OUT_2_port, data_out(1) => 
                           ALU_OUTPUT_OUT_1_port, data_out(0) => 
                           ALU_OUTPUT_OUT_0_port);
   NPC3 : gen_reg_N32_2 port map( clk => CLK, rst => RST, ld => MEM_OUTREG_EN, 
                           data_in(31) => NPC_IN(31), data_in(30) => NPC_IN(30)
                           , data_in(29) => NPC_IN(29), data_in(28) => 
                           NPC_IN(28), data_in(27) => NPC_IN(27), data_in(26) 
                           => NPC_IN(26), data_in(25) => NPC_IN(25), 
                           data_in(24) => NPC_IN(24), data_in(23) => NPC_IN(23)
                           , data_in(22) => NPC_IN(22), data_in(21) => 
                           NPC_IN(21), data_in(20) => NPC_IN(20), data_in(19) 
                           => NPC_IN(19), data_in(18) => NPC_IN(18), 
                           data_in(17) => NPC_IN(17), data_in(16) => NPC_IN(16)
                           , data_in(15) => NPC_IN(15), data_in(14) => 
                           NPC_IN(14), data_in(13) => NPC_IN(13), data_in(12) 
                           => NPC_IN(12), data_in(11) => NPC_IN(11), 
                           data_in(10) => NPC_IN(10), data_in(9) => NPC_IN(9), 
                           data_in(8) => NPC_IN(8), data_in(7) => NPC_IN(7), 
                           data_in(6) => NPC_IN(6), data_in(5) => NPC_IN(5), 
                           data_in(4) => NPC_IN(4), data_in(3) => NPC_IN(3), 
                           data_in(2) => NPC_IN(2), data_in(1) => NPC_IN(1), 
                           data_in(0) => NPC_IN(0), data_out(31) => NPC_OUT(31)
                           , data_out(30) => NPC_OUT(30), data_out(29) => 
                           NPC_OUT(29), data_out(28) => NPC_OUT(28), 
                           data_out(27) => NPC_OUT(27), data_out(26) => 
                           NPC_OUT(26), data_out(25) => NPC_OUT(25), 
                           data_out(24) => NPC_OUT(24), data_out(23) => 
                           NPC_OUT(23), data_out(22) => NPC_OUT(22), 
                           data_out(21) => NPC_OUT(21), data_out(20) => 
                           NPC_OUT(20), data_out(19) => NPC_OUT(19), 
                           data_out(18) => NPC_OUT(18), data_out(17) => 
                           NPC_OUT(17), data_out(16) => NPC_OUT(16), 
                           data_out(15) => NPC_OUT(15), data_out(14) => 
                           NPC_OUT(14), data_out(13) => NPC_OUT(13), 
                           data_out(12) => NPC_OUT(12), data_out(11) => 
                           NPC_OUT(11), data_out(10) => NPC_OUT(10), 
                           data_out(9) => NPC_OUT(9), data_out(8) => NPC_OUT(8)
                           , data_out(7) => NPC_OUT(7), data_out(6) => 
                           NPC_OUT(6), data_out(5) => NPC_OUT(5), data_out(4) 
                           => NPC_OUT(4), data_out(3) => NPC_OUT(3), 
                           data_out(2) => NPC_OUT(2), data_out(1) => NPC_OUT(1)
                           , data_out(0) => NPC_OUT(0));
   IR3 : gen_reg_N5_2 port map( clk => CLK, rst => RST, ld => MEM_OUTREG_EN, 
                           data_in(4) => IR_IN(4), data_in(3) => IR_IN(3), 
                           data_in(2) => IR_IN(2), data_in(1) => IR_IN(1), 
                           data_in(0) => IR_IN(0), data_out(4) => IR_OUT(4), 
                           data_out(3) => IR_OUT(3), data_out(2) => IR_OUT(2), 
                           data_out(1) => IR_OUT(1), data_out(0) => IR_OUT(0));
   SIGN_EXT_BLOCK : sign_ext_alt_N_IN016_N_IN18_N_OUT32 port map( ctrl_in => 
                           BYTE_LEN_IN(0), zero_padding => ZERO_PADDING4, 
                           data_in(15) => MEM_DATA_OUT_INT(15), data_in(14) => 
                           MEM_DATA_OUT_INT(14), data_in(13) => 
                           MEM_DATA_OUT_INT(13), data_in(12) => 
                           MEM_DATA_OUT_INT(12), data_in(11) => 
                           MEM_DATA_OUT_INT(11), data_in(10) => 
                           MEM_DATA_OUT_INT(10), data_in(9) => 
                           MEM_DATA_OUT_INT(9), data_in(8) => 
                           MEM_DATA_OUT_INT(8), data_in(7) => 
                           MEM_DATA_OUT_INT(7), data_in(6) => 
                           MEM_DATA_OUT_INT(6), data_in(5) => 
                           MEM_DATA_OUT_INT(5), data_in(4) => 
                           MEM_DATA_OUT_INT(4), data_in(3) => 
                           MEM_DATA_OUT_INT(3), data_in(2) => 
                           MEM_DATA_OUT_INT(2), data_in(1) => 
                           MEM_DATA_OUT_INT(1), data_in(0) => 
                           MEM_DATA_OUT_INT(0), data_ext(31) => 
                           SIGN_EXT_OUT_31_port, data_ext(30) => 
                           SIGN_EXT_OUT_30_port, data_ext(29) => 
                           SIGN_EXT_OUT_29_port, data_ext(28) => 
                           SIGN_EXT_OUT_28_port, data_ext(27) => 
                           SIGN_EXT_OUT_27_port, data_ext(26) => 
                           SIGN_EXT_OUT_26_port, data_ext(25) => 
                           SIGN_EXT_OUT_25_port, data_ext(24) => 
                           SIGN_EXT_OUT_24_port, data_ext(23) => 
                           SIGN_EXT_OUT_23_port, data_ext(22) => 
                           SIGN_EXT_OUT_22_port, data_ext(21) => 
                           SIGN_EXT_OUT_21_port, data_ext(20) => 
                           SIGN_EXT_OUT_20_port, data_ext(19) => 
                           SIGN_EXT_OUT_19_port, data_ext(18) => 
                           SIGN_EXT_OUT_18_port, data_ext(17) => 
                           SIGN_EXT_OUT_17_port, data_ext(16) => 
                           SIGN_EXT_OUT_16_port, data_ext(15) => 
                           SIGN_EXT_OUT_15_port, data_ext(14) => 
                           SIGN_EXT_OUT_14_port, data_ext(13) => 
                           SIGN_EXT_OUT_13_port, data_ext(12) => 
                           SIGN_EXT_OUT_12_port, data_ext(11) => 
                           SIGN_EXT_OUT_11_port, data_ext(10) => 
                           SIGN_EXT_OUT_10_port, data_ext(9) => 
                           SIGN_EXT_OUT_9_port, data_ext(8) => 
                           SIGN_EXT_OUT_8_port, data_ext(7) => 
                           SIGN_EXT_OUT_7_port, data_ext(6) => 
                           SIGN_EXT_OUT_6_port, data_ext(5) => 
                           SIGN_EXT_OUT_5_port, data_ext(4) => 
                           SIGN_EXT_OUT_4_port, data_ext(3) => 
                           SIGN_EXT_OUT_3_port, data_ext(2) => 
                           SIGN_EXT_OUT_2_port, data_ext(1) => 
                           SIGN_EXT_OUT_1_port, data_ext(0) => 
                           SIGN_EXT_OUT_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity EXE_STAGE_N_BITS_DATA32_RF_ADDR5 is

   port( CLK, RST, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN : in 
         std_logic;  ALU_OPCODE : in std_logic_vector (0 to 6);  NPC2_IN, 
         NPC1_MUXA_IN, REGA_MUXA_IN, REGB_MUXB_IN, IMM_MUXB_IN, PAD_IN : in 
         std_logic_vector (31 downto 0);  IR2_IN : in std_logic_vector (4 
         downto 0);  NPC2_OUT : out std_logic_vector (31 downto 0);  
         ZERO_OP_OUT : out std_logic;  ALU_OUT, PAD_OUT : out std_logic_vector 
         (31 downto 0);  IR2_OUT : out std_logic_vector (4 downto 0);  N_FLAG, 
         Z_FLAG, C_FLAG, V_FLAG : out std_logic);

end EXE_STAGE_N_BITS_DATA32_RF_ADDR5;

architecture SYN_STRUCTURAL of EXE_STAGE_N_BITS_DATA32_RF_ADDR5 is

   component gen_reg_N5_3
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 
            downto 0);  data_out : out std_logic_vector (4 downto 0));
   end component;
   
   component gen_reg_N32_4
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component cpsr
      port( clk, rst, ld, FL3, FL2, FL1, FL0 : in std_logic;  N, Z, C, V : out 
            std_logic);
   end component;
   
   component gen_reg_N32_5
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_N32
      port( ALU_OPCODE : in std_logic_vector (0 to 6);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  NEG, ZERO, CARRY, OVF : out 
            std_logic;  OUTALU : out std_logic_vector (31 downto 0));
   end component;
   
   component gen_mux21_N32_3
      port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m :
            out std_logic_vector (31 downto 0));
   end component;
   
   component gen_mux21_N32_0
      port( sel : in std_logic;  x, y : in std_logic_vector (31 downto 0);  m :
            out std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N1_0
      port( clk, rst, ld, data_in : in std_logic;  data_out : out std_logic);
   end component;
   
   component cond_branch
      port( cond_in, jump_in, ctrl_in : in std_logic;  ctrl_out : out std_logic
            );
   end component;
   
   component zero_check_N32
      port( data_in : in std_logic_vector (31 downto 0);  ctrl_out : out 
            std_logic);
   end component;
   
   component gen_reg_N32_6
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal BRANCH_TAKEN, ZERO_REG_IN_0_port, MUXA_OUT_INT_31_port, 
      MUXA_OUT_INT_30_port, MUXA_OUT_INT_29_port, MUXA_OUT_INT_28_port, 
      MUXA_OUT_INT_27_port, MUXA_OUT_INT_26_port, MUXA_OUT_INT_25_port, 
      MUXA_OUT_INT_24_port, MUXA_OUT_INT_23_port, MUXA_OUT_INT_22_port, 
      MUXA_OUT_INT_21_port, MUXA_OUT_INT_20_port, MUXA_OUT_INT_19_port, 
      MUXA_OUT_INT_18_port, MUXA_OUT_INT_17_port, MUXA_OUT_INT_16_port, 
      MUXA_OUT_INT_15_port, MUXA_OUT_INT_14_port, MUXA_OUT_INT_13_port, 
      MUXA_OUT_INT_12_port, MUXA_OUT_INT_11_port, MUXA_OUT_INT_10_port, 
      MUXA_OUT_INT_9_port, MUXA_OUT_INT_8_port, MUXA_OUT_INT_7_port, 
      MUXA_OUT_INT_6_port, MUXA_OUT_INT_5_port, MUXA_OUT_INT_4_port, 
      MUXA_OUT_INT_3_port, MUXA_OUT_INT_2_port, MUXA_OUT_INT_1_port, 
      MUXA_OUT_INT_0_port, MUXB_OUT_INT_31_port, MUXB_OUT_INT_30_port, 
      MUXB_OUT_INT_29_port, MUXB_OUT_INT_28_port, MUXB_OUT_INT_27_port, 
      MUXB_OUT_INT_26_port, MUXB_OUT_INT_25_port, MUXB_OUT_INT_24_port, 
      MUXB_OUT_INT_23_port, MUXB_OUT_INT_22_port, MUXB_OUT_INT_21_port, 
      MUXB_OUT_INT_20_port, MUXB_OUT_INT_19_port, MUXB_OUT_INT_18_port, 
      MUXB_OUT_INT_17_port, MUXB_OUT_INT_16_port, MUXB_OUT_INT_15_port, 
      MUXB_OUT_INT_14_port, MUXB_OUT_INT_13_port, MUXB_OUT_INT_12_port, 
      MUXB_OUT_INT_11_port, MUXB_OUT_INT_10_port, MUXB_OUT_INT_9_port, 
      MUXB_OUT_INT_8_port, MUXB_OUT_INT_7_port, MUXB_OUT_INT_6_port, 
      MUXB_OUT_INT_5_port, MUXB_OUT_INT_4_port, MUXB_OUT_INT_3_port, 
      MUXB_OUT_INT_2_port, MUXB_OUT_INT_1_port, MUXB_OUT_INT_0_port, NEG_INT, 
      ZERO_INT, CARRY_INT, OVF_INT, ALU_OUT_INT_31_port, ALU_OUT_INT_30_port, 
      ALU_OUT_INT_29_port, ALU_OUT_INT_28_port, ALU_OUT_INT_27_port, 
      ALU_OUT_INT_26_port, ALU_OUT_INT_25_port, ALU_OUT_INT_24_port, 
      ALU_OUT_INT_23_port, ALU_OUT_INT_22_port, ALU_OUT_INT_21_port, 
      ALU_OUT_INT_20_port, ALU_OUT_INT_19_port, ALU_OUT_INT_18_port, 
      ALU_OUT_INT_17_port, ALU_OUT_INT_16_port, ALU_OUT_INT_15_port, 
      ALU_OUT_INT_14_port, ALU_OUT_INT_13_port, ALU_OUT_INT_12_port, 
      ALU_OUT_INT_11_port, ALU_OUT_INT_10_port, ALU_OUT_INT_9_port, 
      ALU_OUT_INT_8_port, ALU_OUT_INT_7_port, ALU_OUT_INT_6_port, 
      ALU_OUT_INT_5_port, ALU_OUT_INT_4_port, ALU_OUT_INT_3_port, 
      ALU_OUT_INT_2_port, ALU_OUT_INT_1_port, ALU_OUT_INT_0_port : std_logic;

begin
   
   NPC2 : gen_reg_N32_6 port map( clk => CLK, rst => RST, ld => EXE_OUTREG_EN, 
                           data_in(31) => NPC2_IN(31), data_in(30) => 
                           NPC2_IN(30), data_in(29) => NPC2_IN(29), data_in(28)
                           => NPC2_IN(28), data_in(27) => NPC2_IN(27), 
                           data_in(26) => NPC2_IN(26), data_in(25) => 
                           NPC2_IN(25), data_in(24) => NPC2_IN(24), data_in(23)
                           => NPC2_IN(23), data_in(22) => NPC2_IN(22), 
                           data_in(21) => NPC2_IN(21), data_in(20) => 
                           NPC2_IN(20), data_in(19) => NPC2_IN(19), data_in(18)
                           => NPC2_IN(18), data_in(17) => NPC2_IN(17), 
                           data_in(16) => NPC2_IN(16), data_in(15) => 
                           NPC2_IN(15), data_in(14) => NPC2_IN(14), data_in(13)
                           => NPC2_IN(13), data_in(12) => NPC2_IN(12), 
                           data_in(11) => NPC2_IN(11), data_in(10) => 
                           NPC2_IN(10), data_in(9) => NPC2_IN(9), data_in(8) =>
                           NPC2_IN(8), data_in(7) => NPC2_IN(7), data_in(6) => 
                           NPC2_IN(6), data_in(5) => NPC2_IN(5), data_in(4) => 
                           NPC2_IN(4), data_in(3) => NPC2_IN(3), data_in(2) => 
                           NPC2_IN(2), data_in(1) => NPC2_IN(1), data_in(0) => 
                           NPC2_IN(0), data_out(31) => NPC2_OUT(31), 
                           data_out(30) => NPC2_OUT(30), data_out(29) => 
                           NPC2_OUT(29), data_out(28) => NPC2_OUT(28), 
                           data_out(27) => NPC2_OUT(27), data_out(26) => 
                           NPC2_OUT(26), data_out(25) => NPC2_OUT(25), 
                           data_out(24) => NPC2_OUT(24), data_out(23) => 
                           NPC2_OUT(23), data_out(22) => NPC2_OUT(22), 
                           data_out(21) => NPC2_OUT(21), data_out(20) => 
                           NPC2_OUT(20), data_out(19) => NPC2_OUT(19), 
                           data_out(18) => NPC2_OUT(18), data_out(17) => 
                           NPC2_OUT(17), data_out(16) => NPC2_OUT(16), 
                           data_out(15) => NPC2_OUT(15), data_out(14) => 
                           NPC2_OUT(14), data_out(13) => NPC2_OUT(13), 
                           data_out(12) => NPC2_OUT(12), data_out(11) => 
                           NPC2_OUT(11), data_out(10) => NPC2_OUT(10), 
                           data_out(9) => NPC2_OUT(9), data_out(8) => 
                           NPC2_OUT(8), data_out(7) => NPC2_OUT(7), data_out(6)
                           => NPC2_OUT(6), data_out(5) => NPC2_OUT(5), 
                           data_out(4) => NPC2_OUT(4), data_out(3) => 
                           NPC2_OUT(3), data_out(2) => NPC2_OUT(2), data_out(1)
                           => NPC2_OUT(1), data_out(0) => NPC2_OUT(0));
   ZERO : zero_check_N32 port map( data_in(31) => REGA_MUXA_IN(31), data_in(30)
                           => REGA_MUXA_IN(30), data_in(29) => REGA_MUXA_IN(29)
                           , data_in(28) => REGA_MUXA_IN(28), data_in(27) => 
                           REGA_MUXA_IN(27), data_in(26) => REGA_MUXA_IN(26), 
                           data_in(25) => REGA_MUXA_IN(25), data_in(24) => 
                           REGA_MUXA_IN(24), data_in(23) => REGA_MUXA_IN(23), 
                           data_in(22) => REGA_MUXA_IN(22), data_in(21) => 
                           REGA_MUXA_IN(21), data_in(20) => REGA_MUXA_IN(20), 
                           data_in(19) => REGA_MUXA_IN(19), data_in(18) => 
                           REGA_MUXA_IN(18), data_in(17) => REGA_MUXA_IN(17), 
                           data_in(16) => REGA_MUXA_IN(16), data_in(15) => 
                           REGA_MUXA_IN(15), data_in(14) => REGA_MUXA_IN(14), 
                           data_in(13) => REGA_MUXA_IN(13), data_in(12) => 
                           REGA_MUXA_IN(12), data_in(11) => REGA_MUXA_IN(11), 
                           data_in(10) => REGA_MUXA_IN(10), data_in(9) => 
                           REGA_MUXA_IN(9), data_in(8) => REGA_MUXA_IN(8), 
                           data_in(7) => REGA_MUXA_IN(7), data_in(6) => 
                           REGA_MUXA_IN(6), data_in(5) => REGA_MUXA_IN(5), 
                           data_in(4) => REGA_MUXA_IN(4), data_in(3) => 
                           REGA_MUXA_IN(3), data_in(2) => REGA_MUXA_IN(2), 
                           data_in(1) => REGA_MUXA_IN(1), data_in(0) => 
                           REGA_MUXA_IN(0), ctrl_out => BRANCH_TAKEN);
   COND : cond_branch port map( cond_in => EQ_COND, jump_in => JUMP_EN, ctrl_in
                           => BRANCH_TAKEN, ctrl_out => ZERO_REG_IN_0_port);
   ZOP : gen_reg_N1_0 port map( clk => CLK, rst => RST, ld => EXE_OUTREG_EN, 
                           data_in => ZERO_REG_IN_0_port, data_out => 
                           ZERO_OP_OUT);
   MUXA : gen_mux21_N32_0 port map( sel => MUXA_SEL, x(31) => NPC1_MUXA_IN(31),
                           x(30) => NPC1_MUXA_IN(30), x(29) => NPC1_MUXA_IN(29)
                           , x(28) => NPC1_MUXA_IN(28), x(27) => 
                           NPC1_MUXA_IN(27), x(26) => NPC1_MUXA_IN(26), x(25) 
                           => NPC1_MUXA_IN(25), x(24) => NPC1_MUXA_IN(24), 
                           x(23) => NPC1_MUXA_IN(23), x(22) => NPC1_MUXA_IN(22)
                           , x(21) => NPC1_MUXA_IN(21), x(20) => 
                           NPC1_MUXA_IN(20), x(19) => NPC1_MUXA_IN(19), x(18) 
                           => NPC1_MUXA_IN(18), x(17) => NPC1_MUXA_IN(17), 
                           x(16) => NPC1_MUXA_IN(16), x(15) => NPC1_MUXA_IN(15)
                           , x(14) => NPC1_MUXA_IN(14), x(13) => 
                           NPC1_MUXA_IN(13), x(12) => NPC1_MUXA_IN(12), x(11) 
                           => NPC1_MUXA_IN(11), x(10) => NPC1_MUXA_IN(10), x(9)
                           => NPC1_MUXA_IN(9), x(8) => NPC1_MUXA_IN(8), x(7) =>
                           NPC1_MUXA_IN(7), x(6) => NPC1_MUXA_IN(6), x(5) => 
                           NPC1_MUXA_IN(5), x(4) => NPC1_MUXA_IN(4), x(3) => 
                           NPC1_MUXA_IN(3), x(2) => NPC1_MUXA_IN(2), x(1) => 
                           NPC1_MUXA_IN(1), x(0) => NPC1_MUXA_IN(0), y(31) => 
                           REGA_MUXA_IN(31), y(30) => REGA_MUXA_IN(30), y(29) 
                           => REGA_MUXA_IN(29), y(28) => REGA_MUXA_IN(28), 
                           y(27) => REGA_MUXA_IN(27), y(26) => REGA_MUXA_IN(26)
                           , y(25) => REGA_MUXA_IN(25), y(24) => 
                           REGA_MUXA_IN(24), y(23) => REGA_MUXA_IN(23), y(22) 
                           => REGA_MUXA_IN(22), y(21) => REGA_MUXA_IN(21), 
                           y(20) => REGA_MUXA_IN(20), y(19) => REGA_MUXA_IN(19)
                           , y(18) => REGA_MUXA_IN(18), y(17) => 
                           REGA_MUXA_IN(17), y(16) => REGA_MUXA_IN(16), y(15) 
                           => REGA_MUXA_IN(15), y(14) => REGA_MUXA_IN(14), 
                           y(13) => REGA_MUXA_IN(13), y(12) => REGA_MUXA_IN(12)
                           , y(11) => REGA_MUXA_IN(11), y(10) => 
                           REGA_MUXA_IN(10), y(9) => REGA_MUXA_IN(9), y(8) => 
                           REGA_MUXA_IN(8), y(7) => REGA_MUXA_IN(7), y(6) => 
                           REGA_MUXA_IN(6), y(5) => REGA_MUXA_IN(5), y(4) => 
                           REGA_MUXA_IN(4), y(3) => REGA_MUXA_IN(3), y(2) => 
                           REGA_MUXA_IN(2), y(1) => REGA_MUXA_IN(1), y(0) => 
                           REGA_MUXA_IN(0), m(31) => MUXA_OUT_INT_31_port, 
                           m(30) => MUXA_OUT_INT_30_port, m(29) => 
                           MUXA_OUT_INT_29_port, m(28) => MUXA_OUT_INT_28_port,
                           m(27) => MUXA_OUT_INT_27_port, m(26) => 
                           MUXA_OUT_INT_26_port, m(25) => MUXA_OUT_INT_25_port,
                           m(24) => MUXA_OUT_INT_24_port, m(23) => 
                           MUXA_OUT_INT_23_port, m(22) => MUXA_OUT_INT_22_port,
                           m(21) => MUXA_OUT_INT_21_port, m(20) => 
                           MUXA_OUT_INT_20_port, m(19) => MUXA_OUT_INT_19_port,
                           m(18) => MUXA_OUT_INT_18_port, m(17) => 
                           MUXA_OUT_INT_17_port, m(16) => MUXA_OUT_INT_16_port,
                           m(15) => MUXA_OUT_INT_15_port, m(14) => 
                           MUXA_OUT_INT_14_port, m(13) => MUXA_OUT_INT_13_port,
                           m(12) => MUXA_OUT_INT_12_port, m(11) => 
                           MUXA_OUT_INT_11_port, m(10) => MUXA_OUT_INT_10_port,
                           m(9) => MUXA_OUT_INT_9_port, m(8) => 
                           MUXA_OUT_INT_8_port, m(7) => MUXA_OUT_INT_7_port, 
                           m(6) => MUXA_OUT_INT_6_port, m(5) => 
                           MUXA_OUT_INT_5_port, m(4) => MUXA_OUT_INT_4_port, 
                           m(3) => MUXA_OUT_INT_3_port, m(2) => 
                           MUXA_OUT_INT_2_port, m(1) => MUXA_OUT_INT_1_port, 
                           m(0) => MUXA_OUT_INT_0_port);
   MUXB : gen_mux21_N32_3 port map( sel => MUXB_SEL, x(31) => REGB_MUXB_IN(31),
                           x(30) => REGB_MUXB_IN(30), x(29) => REGB_MUXB_IN(29)
                           , x(28) => REGB_MUXB_IN(28), x(27) => 
                           REGB_MUXB_IN(27), x(26) => REGB_MUXB_IN(26), x(25) 
                           => REGB_MUXB_IN(25), x(24) => REGB_MUXB_IN(24), 
                           x(23) => REGB_MUXB_IN(23), x(22) => REGB_MUXB_IN(22)
                           , x(21) => REGB_MUXB_IN(21), x(20) => 
                           REGB_MUXB_IN(20), x(19) => REGB_MUXB_IN(19), x(18) 
                           => REGB_MUXB_IN(18), x(17) => REGB_MUXB_IN(17), 
                           x(16) => REGB_MUXB_IN(16), x(15) => REGB_MUXB_IN(15)
                           , x(14) => REGB_MUXB_IN(14), x(13) => 
                           REGB_MUXB_IN(13), x(12) => REGB_MUXB_IN(12), x(11) 
                           => REGB_MUXB_IN(11), x(10) => REGB_MUXB_IN(10), x(9)
                           => REGB_MUXB_IN(9), x(8) => REGB_MUXB_IN(8), x(7) =>
                           REGB_MUXB_IN(7), x(6) => REGB_MUXB_IN(6), x(5) => 
                           REGB_MUXB_IN(5), x(4) => REGB_MUXB_IN(4), x(3) => 
                           REGB_MUXB_IN(3), x(2) => REGB_MUXB_IN(2), x(1) => 
                           REGB_MUXB_IN(1), x(0) => REGB_MUXB_IN(0), y(31) => 
                           IMM_MUXB_IN(31), y(30) => IMM_MUXB_IN(30), y(29) => 
                           IMM_MUXB_IN(29), y(28) => IMM_MUXB_IN(28), y(27) => 
                           IMM_MUXB_IN(27), y(26) => IMM_MUXB_IN(26), y(25) => 
                           IMM_MUXB_IN(25), y(24) => IMM_MUXB_IN(24), y(23) => 
                           IMM_MUXB_IN(23), y(22) => IMM_MUXB_IN(22), y(21) => 
                           IMM_MUXB_IN(21), y(20) => IMM_MUXB_IN(20), y(19) => 
                           IMM_MUXB_IN(19), y(18) => IMM_MUXB_IN(18), y(17) => 
                           IMM_MUXB_IN(17), y(16) => IMM_MUXB_IN(16), y(15) => 
                           IMM_MUXB_IN(15), y(14) => IMM_MUXB_IN(14), y(13) => 
                           IMM_MUXB_IN(13), y(12) => IMM_MUXB_IN(12), y(11) => 
                           IMM_MUXB_IN(11), y(10) => IMM_MUXB_IN(10), y(9) => 
                           IMM_MUXB_IN(9), y(8) => IMM_MUXB_IN(8), y(7) => 
                           IMM_MUXB_IN(7), y(6) => IMM_MUXB_IN(6), y(5) => 
                           IMM_MUXB_IN(5), y(4) => IMM_MUXB_IN(4), y(3) => 
                           IMM_MUXB_IN(3), y(2) => IMM_MUXB_IN(2), y(1) => 
                           IMM_MUXB_IN(1), y(0) => IMM_MUXB_IN(0), m(31) => 
                           MUXB_OUT_INT_31_port, m(30) => MUXB_OUT_INT_30_port,
                           m(29) => MUXB_OUT_INT_29_port, m(28) => 
                           MUXB_OUT_INT_28_port, m(27) => MUXB_OUT_INT_27_port,
                           m(26) => MUXB_OUT_INT_26_port, m(25) => 
                           MUXB_OUT_INT_25_port, m(24) => MUXB_OUT_INT_24_port,
                           m(23) => MUXB_OUT_INT_23_port, m(22) => 
                           MUXB_OUT_INT_22_port, m(21) => MUXB_OUT_INT_21_port,
                           m(20) => MUXB_OUT_INT_20_port, m(19) => 
                           MUXB_OUT_INT_19_port, m(18) => MUXB_OUT_INT_18_port,
                           m(17) => MUXB_OUT_INT_17_port, m(16) => 
                           MUXB_OUT_INT_16_port, m(15) => MUXB_OUT_INT_15_port,
                           m(14) => MUXB_OUT_INT_14_port, m(13) => 
                           MUXB_OUT_INT_13_port, m(12) => MUXB_OUT_INT_12_port,
                           m(11) => MUXB_OUT_INT_11_port, m(10) => 
                           MUXB_OUT_INT_10_port, m(9) => MUXB_OUT_INT_9_port, 
                           m(8) => MUXB_OUT_INT_8_port, m(7) => 
                           MUXB_OUT_INT_7_port, m(6) => MUXB_OUT_INT_6_port, 
                           m(5) => MUXB_OUT_INT_5_port, m(4) => 
                           MUXB_OUT_INT_4_port, m(3) => MUXB_OUT_INT_3_port, 
                           m(2) => MUXB_OUT_INT_2_port, m(1) => 
                           MUXB_OUT_INT_1_port, m(0) => MUXB_OUT_INT_0_port);
   ALRITH_LOG_U : ALU_N32 port map( ALU_OPCODE(0) => ALU_OPCODE(0), 
                           ALU_OPCODE(1) => ALU_OPCODE(1), ALU_OPCODE(2) => 
                           ALU_OPCODE(2), ALU_OPCODE(3) => ALU_OPCODE(3), 
                           ALU_OPCODE(4) => ALU_OPCODE(4), ALU_OPCODE(5) => 
                           ALU_OPCODE(5), ALU_OPCODE(6) => ALU_OPCODE(6), 
                           DATA1(31) => MUXA_OUT_INT_31_port, DATA1(30) => 
                           MUXA_OUT_INT_30_port, DATA1(29) => 
                           MUXA_OUT_INT_29_port, DATA1(28) => 
                           MUXA_OUT_INT_28_port, DATA1(27) => 
                           MUXA_OUT_INT_27_port, DATA1(26) => 
                           MUXA_OUT_INT_26_port, DATA1(25) => 
                           MUXA_OUT_INT_25_port, DATA1(24) => 
                           MUXA_OUT_INT_24_port, DATA1(23) => 
                           MUXA_OUT_INT_23_port, DATA1(22) => 
                           MUXA_OUT_INT_22_port, DATA1(21) => 
                           MUXA_OUT_INT_21_port, DATA1(20) => 
                           MUXA_OUT_INT_20_port, DATA1(19) => 
                           MUXA_OUT_INT_19_port, DATA1(18) => 
                           MUXA_OUT_INT_18_port, DATA1(17) => 
                           MUXA_OUT_INT_17_port, DATA1(16) => 
                           MUXA_OUT_INT_16_port, DATA1(15) => 
                           MUXA_OUT_INT_15_port, DATA1(14) => 
                           MUXA_OUT_INT_14_port, DATA1(13) => 
                           MUXA_OUT_INT_13_port, DATA1(12) => 
                           MUXA_OUT_INT_12_port, DATA1(11) => 
                           MUXA_OUT_INT_11_port, DATA1(10) => 
                           MUXA_OUT_INT_10_port, DATA1(9) => 
                           MUXA_OUT_INT_9_port, DATA1(8) => MUXA_OUT_INT_8_port
                           , DATA1(7) => MUXA_OUT_INT_7_port, DATA1(6) => 
                           MUXA_OUT_INT_6_port, DATA1(5) => MUXA_OUT_INT_5_port
                           , DATA1(4) => MUXA_OUT_INT_4_port, DATA1(3) => 
                           MUXA_OUT_INT_3_port, DATA1(2) => MUXA_OUT_INT_2_port
                           , DATA1(1) => MUXA_OUT_INT_1_port, DATA1(0) => 
                           MUXA_OUT_INT_0_port, DATA2(31) => 
                           MUXB_OUT_INT_31_port, DATA2(30) => 
                           MUXB_OUT_INT_30_port, DATA2(29) => 
                           MUXB_OUT_INT_29_port, DATA2(28) => 
                           MUXB_OUT_INT_28_port, DATA2(27) => 
                           MUXB_OUT_INT_27_port, DATA2(26) => 
                           MUXB_OUT_INT_26_port, DATA2(25) => 
                           MUXB_OUT_INT_25_port, DATA2(24) => 
                           MUXB_OUT_INT_24_port, DATA2(23) => 
                           MUXB_OUT_INT_23_port, DATA2(22) => 
                           MUXB_OUT_INT_22_port, DATA2(21) => 
                           MUXB_OUT_INT_21_port, DATA2(20) => 
                           MUXB_OUT_INT_20_port, DATA2(19) => 
                           MUXB_OUT_INT_19_port, DATA2(18) => 
                           MUXB_OUT_INT_18_port, DATA2(17) => 
                           MUXB_OUT_INT_17_port, DATA2(16) => 
                           MUXB_OUT_INT_16_port, DATA2(15) => 
                           MUXB_OUT_INT_15_port, DATA2(14) => 
                           MUXB_OUT_INT_14_port, DATA2(13) => 
                           MUXB_OUT_INT_13_port, DATA2(12) => 
                           MUXB_OUT_INT_12_port, DATA2(11) => 
                           MUXB_OUT_INT_11_port, DATA2(10) => 
                           MUXB_OUT_INT_10_port, DATA2(9) => 
                           MUXB_OUT_INT_9_port, DATA2(8) => MUXB_OUT_INT_8_port
                           , DATA2(7) => MUXB_OUT_INT_7_port, DATA2(6) => 
                           MUXB_OUT_INT_6_port, DATA2(5) => MUXB_OUT_INT_5_port
                           , DATA2(4) => MUXB_OUT_INT_4_port, DATA2(3) => 
                           MUXB_OUT_INT_3_port, DATA2(2) => MUXB_OUT_INT_2_port
                           , DATA2(1) => MUXB_OUT_INT_1_port, DATA2(0) => 
                           MUXB_OUT_INT_0_port, NEG => NEG_INT, ZERO => 
                           ZERO_INT, CARRY => CARRY_INT, OVF => OVF_INT, 
                           OUTALU(31) => ALU_OUT_INT_31_port, OUTALU(30) => 
                           ALU_OUT_INT_30_port, OUTALU(29) => 
                           ALU_OUT_INT_29_port, OUTALU(28) => 
                           ALU_OUT_INT_28_port, OUTALU(27) => 
                           ALU_OUT_INT_27_port, OUTALU(26) => 
                           ALU_OUT_INT_26_port, OUTALU(25) => 
                           ALU_OUT_INT_25_port, OUTALU(24) => 
                           ALU_OUT_INT_24_port, OUTALU(23) => 
                           ALU_OUT_INT_23_port, OUTALU(22) => 
                           ALU_OUT_INT_22_port, OUTALU(21) => 
                           ALU_OUT_INT_21_port, OUTALU(20) => 
                           ALU_OUT_INT_20_port, OUTALU(19) => 
                           ALU_OUT_INT_19_port, OUTALU(18) => 
                           ALU_OUT_INT_18_port, OUTALU(17) => 
                           ALU_OUT_INT_17_port, OUTALU(16) => 
                           ALU_OUT_INT_16_port, OUTALU(15) => 
                           ALU_OUT_INT_15_port, OUTALU(14) => 
                           ALU_OUT_INT_14_port, OUTALU(13) => 
                           ALU_OUT_INT_13_port, OUTALU(12) => 
                           ALU_OUT_INT_12_port, OUTALU(11) => 
                           ALU_OUT_INT_11_port, OUTALU(10) => 
                           ALU_OUT_INT_10_port, OUTALU(9) => ALU_OUT_INT_9_port
                           , OUTALU(8) => ALU_OUT_INT_8_port, OUTALU(7) => 
                           ALU_OUT_INT_7_port, OUTALU(6) => ALU_OUT_INT_6_port,
                           OUTALU(5) => ALU_OUT_INT_5_port, OUTALU(4) => 
                           ALU_OUT_INT_4_port, OUTALU(3) => ALU_OUT_INT_3_port,
                           OUTALU(2) => ALU_OUT_INT_2_port, OUTALU(1) => 
                           ALU_OUT_INT_1_port, OUTALU(0) => ALU_OUT_INT_0_port)
                           ;
   ALU_OUTPUT : gen_reg_N32_5 port map( clk => CLK, rst => RST, ld => 
                           EXE_OUTREG_EN, data_in(31) => ALU_OUT_INT_31_port, 
                           data_in(30) => ALU_OUT_INT_30_port, data_in(29) => 
                           ALU_OUT_INT_29_port, data_in(28) => 
                           ALU_OUT_INT_28_port, data_in(27) => 
                           ALU_OUT_INT_27_port, data_in(26) => 
                           ALU_OUT_INT_26_port, data_in(25) => 
                           ALU_OUT_INT_25_port, data_in(24) => 
                           ALU_OUT_INT_24_port, data_in(23) => 
                           ALU_OUT_INT_23_port, data_in(22) => 
                           ALU_OUT_INT_22_port, data_in(21) => 
                           ALU_OUT_INT_21_port, data_in(20) => 
                           ALU_OUT_INT_20_port, data_in(19) => 
                           ALU_OUT_INT_19_port, data_in(18) => 
                           ALU_OUT_INT_18_port, data_in(17) => 
                           ALU_OUT_INT_17_port, data_in(16) => 
                           ALU_OUT_INT_16_port, data_in(15) => 
                           ALU_OUT_INT_15_port, data_in(14) => 
                           ALU_OUT_INT_14_port, data_in(13) => 
                           ALU_OUT_INT_13_port, data_in(12) => 
                           ALU_OUT_INT_12_port, data_in(11) => 
                           ALU_OUT_INT_11_port, data_in(10) => 
                           ALU_OUT_INT_10_port, data_in(9) => 
                           ALU_OUT_INT_9_port, data_in(8) => ALU_OUT_INT_8_port
                           , data_in(7) => ALU_OUT_INT_7_port, data_in(6) => 
                           ALU_OUT_INT_6_port, data_in(5) => ALU_OUT_INT_5_port
                           , data_in(4) => ALU_OUT_INT_4_port, data_in(3) => 
                           ALU_OUT_INT_3_port, data_in(2) => ALU_OUT_INT_2_port
                           , data_in(1) => ALU_OUT_INT_1_port, data_in(0) => 
                           ALU_OUT_INT_0_port, data_out(31) => ALU_OUT(31), 
                           data_out(30) => ALU_OUT(30), data_out(29) => 
                           ALU_OUT(29), data_out(28) => ALU_OUT(28), 
                           data_out(27) => ALU_OUT(27), data_out(26) => 
                           ALU_OUT(26), data_out(25) => ALU_OUT(25), 
                           data_out(24) => ALU_OUT(24), data_out(23) => 
                           ALU_OUT(23), data_out(22) => ALU_OUT(22), 
                           data_out(21) => ALU_OUT(21), data_out(20) => 
                           ALU_OUT(20), data_out(19) => ALU_OUT(19), 
                           data_out(18) => ALU_OUT(18), data_out(17) => 
                           ALU_OUT(17), data_out(16) => ALU_OUT(16), 
                           data_out(15) => ALU_OUT(15), data_out(14) => 
                           ALU_OUT(14), data_out(13) => ALU_OUT(13), 
                           data_out(12) => ALU_OUT(12), data_out(11) => 
                           ALU_OUT(11), data_out(10) => ALU_OUT(10), 
                           data_out(9) => ALU_OUT(9), data_out(8) => ALU_OUT(8)
                           , data_out(7) => ALU_OUT(7), data_out(6) => 
                           ALU_OUT(6), data_out(5) => ALU_OUT(5), data_out(4) 
                           => ALU_OUT(4), data_out(3) => ALU_OUT(3), 
                           data_out(2) => ALU_OUT(2), data_out(1) => ALU_OUT(1)
                           , data_out(0) => ALU_OUT(0));
   ALU_FLAGS : cpsr port map( clk => CLK, rst => RST, ld => EXE_OUTREG_EN, FL3 
                           => NEG_INT, FL2 => ZERO_INT, FL1 => CARRY_INT, FL0 
                           => OVF_INT, N => N_FLAG, Z => Z_FLAG, C => C_FLAG, V
                           => V_FLAG);
   PAD : gen_reg_N32_4 port map( clk => CLK, rst => RST, ld => EXE_OUTREG_EN, 
                           data_in(31) => PAD_IN(31), data_in(30) => PAD_IN(30)
                           , data_in(29) => PAD_IN(29), data_in(28) => 
                           PAD_IN(28), data_in(27) => PAD_IN(27), data_in(26) 
                           => PAD_IN(26), data_in(25) => PAD_IN(25), 
                           data_in(24) => PAD_IN(24), data_in(23) => PAD_IN(23)
                           , data_in(22) => PAD_IN(22), data_in(21) => 
                           PAD_IN(21), data_in(20) => PAD_IN(20), data_in(19) 
                           => PAD_IN(19), data_in(18) => PAD_IN(18), 
                           data_in(17) => PAD_IN(17), data_in(16) => PAD_IN(16)
                           , data_in(15) => PAD_IN(15), data_in(14) => 
                           PAD_IN(14), data_in(13) => PAD_IN(13), data_in(12) 
                           => PAD_IN(12), data_in(11) => PAD_IN(11), 
                           data_in(10) => PAD_IN(10), data_in(9) => PAD_IN(9), 
                           data_in(8) => PAD_IN(8), data_in(7) => PAD_IN(7), 
                           data_in(6) => PAD_IN(6), data_in(5) => PAD_IN(5), 
                           data_in(4) => PAD_IN(4), data_in(3) => PAD_IN(3), 
                           data_in(2) => PAD_IN(2), data_in(1) => PAD_IN(1), 
                           data_in(0) => PAD_IN(0), data_out(31) => PAD_OUT(31)
                           , data_out(30) => PAD_OUT(30), data_out(29) => 
                           PAD_OUT(29), data_out(28) => PAD_OUT(28), 
                           data_out(27) => PAD_OUT(27), data_out(26) => 
                           PAD_OUT(26), data_out(25) => PAD_OUT(25), 
                           data_out(24) => PAD_OUT(24), data_out(23) => 
                           PAD_OUT(23), data_out(22) => PAD_OUT(22), 
                           data_out(21) => PAD_OUT(21), data_out(20) => 
                           PAD_OUT(20), data_out(19) => PAD_OUT(19), 
                           data_out(18) => PAD_OUT(18), data_out(17) => 
                           PAD_OUT(17), data_out(16) => PAD_OUT(16), 
                           data_out(15) => PAD_OUT(15), data_out(14) => 
                           PAD_OUT(14), data_out(13) => PAD_OUT(13), 
                           data_out(12) => PAD_OUT(12), data_out(11) => 
                           PAD_OUT(11), data_out(10) => PAD_OUT(10), 
                           data_out(9) => PAD_OUT(9), data_out(8) => PAD_OUT(8)
                           , data_out(7) => PAD_OUT(7), data_out(6) => 
                           PAD_OUT(6), data_out(5) => PAD_OUT(5), data_out(4) 
                           => PAD_OUT(4), data_out(3) => PAD_OUT(3), 
                           data_out(2) => PAD_OUT(2), data_out(1) => PAD_OUT(1)
                           , data_out(0) => PAD_OUT(0));
   IR2 : gen_reg_N5_3 port map( clk => CLK, rst => RST, ld => EXE_OUTREG_EN, 
                           data_in(4) => IR2_IN(4), data_in(3) => IR2_IN(3), 
                           data_in(2) => IR2_IN(2), data_in(1) => IR2_IN(1), 
                           data_in(0) => IR2_IN(0), data_out(4) => IR2_OUT(4), 
                           data_out(3) => IR2_OUT(3), data_out(2) => IR2_OUT(2)
                           , data_out(1) => IR2_OUT(1), data_out(0) => 
                           IR2_OUT(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16
   is

   port( CLK, RST, JAL_MUX_SEL, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, WR_EN
         , ZERO_PADDING2 : in std_logic;  I_CODE, NPC1_IN, DATA_IN : in 
         std_logic_vector (31 downto 0);  WR_ADDR_IN : in std_logic_vector (4 
         downto 0);  REGA_OUT, REGB_OUT, REGIMM_OUT : out std_logic_vector (31 
         downto 0);  WR_ADDR_OUT : out std_logic_vector (4 downto 0);  NPC1_OUT
         : out std_logic_vector (31 downto 0));

end ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16;

architecture SYN_STRUCTURAL of 
   ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 is

   component gen_mux21_N5
      port( sel : in std_logic;  x, y : in std_logic_vector (4 downto 0);  m : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component sign_ext_N_IN026_N_IN116_N_OUT32
      port( ctrl_in, zero_padding : in std_logic;  data_in : in 
            std_logic_vector (25 downto 0);  data_ext : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component reg_file_Dbits32_Abits5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component gen_reg_N5_0
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (4 
            downto 0);  data_out : out std_logic_vector (4 downto 0));
   end component;
   
   component gen_reg_N32_7
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N32_8
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SIGN_EXT_OUT_31_port, SIGN_EXT_OUT_30_port, SIGN_EXT_OUT_29_port, 
      SIGN_EXT_OUT_28_port, SIGN_EXT_OUT_27_port, SIGN_EXT_OUT_26_port, 
      SIGN_EXT_OUT_25_port, SIGN_EXT_OUT_24_port, SIGN_EXT_OUT_23_port, 
      SIGN_EXT_OUT_22_port, SIGN_EXT_OUT_21_port, SIGN_EXT_OUT_20_port, 
      SIGN_EXT_OUT_19_port, SIGN_EXT_OUT_18_port, SIGN_EXT_OUT_17_port, 
      SIGN_EXT_OUT_16_port, SIGN_EXT_OUT_15_port, SIGN_EXT_OUT_14_port, 
      SIGN_EXT_OUT_13_port, SIGN_EXT_OUT_12_port, SIGN_EXT_OUT_11_port, 
      SIGN_EXT_OUT_10_port, SIGN_EXT_OUT_9_port, SIGN_EXT_OUT_8_port, 
      SIGN_EXT_OUT_7_port, SIGN_EXT_OUT_6_port, SIGN_EXT_OUT_5_port, 
      SIGN_EXT_OUT_4_port, SIGN_EXT_OUT_3_port, SIGN_EXT_OUT_2_port, 
      SIGN_EXT_OUT_1_port, SIGN_EXT_OUT_0_port, MUX_OUT_4_port, MUX_OUT_3_port,
      MUX_OUT_2_port, MUX_OUT_1_port, MUX_OUT_0_port, ADD_WR_4_port, 
      ADD_WR_3_port, ADD_WR_2_port, ADD_WR_1_port, ADD_WR_0_port : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => JAL_MUX_SEL, A2 => WR_ADDR_IN(4), ZN => 
                           ADD_WR_4_port);
   U2 : OR2_X1 port map( A1 => JAL_MUX_SEL, A2 => WR_ADDR_IN(3), ZN => 
                           ADD_WR_3_port);
   U3 : OR2_X1 port map( A1 => JAL_MUX_SEL, A2 => WR_ADDR_IN(2), ZN => 
                           ADD_WR_2_port);
   U4 : OR2_X1 port map( A1 => JAL_MUX_SEL, A2 => WR_ADDR_IN(1), ZN => 
                           ADD_WR_1_port);
   U5 : OR2_X1 port map( A1 => JAL_MUX_SEL, A2 => WR_ADDR_IN(0), ZN => 
                           ADD_WR_0_port);
   NPC1 : gen_reg_N32_8 port map( clk => CLK, rst => RST, ld => DEC_OUTREG_EN, 
                           data_in(31) => NPC1_IN(31), data_in(30) => 
                           NPC1_IN(30), data_in(29) => NPC1_IN(29), data_in(28)
                           => NPC1_IN(28), data_in(27) => NPC1_IN(27), 
                           data_in(26) => NPC1_IN(26), data_in(25) => 
                           NPC1_IN(25), data_in(24) => NPC1_IN(24), data_in(23)
                           => NPC1_IN(23), data_in(22) => NPC1_IN(22), 
                           data_in(21) => NPC1_IN(21), data_in(20) => 
                           NPC1_IN(20), data_in(19) => NPC1_IN(19), data_in(18)
                           => NPC1_IN(18), data_in(17) => NPC1_IN(17), 
                           data_in(16) => NPC1_IN(16), data_in(15) => 
                           NPC1_IN(15), data_in(14) => NPC1_IN(14), data_in(13)
                           => NPC1_IN(13), data_in(12) => NPC1_IN(12), 
                           data_in(11) => NPC1_IN(11), data_in(10) => 
                           NPC1_IN(10), data_in(9) => NPC1_IN(9), data_in(8) =>
                           NPC1_IN(8), data_in(7) => NPC1_IN(7), data_in(6) => 
                           NPC1_IN(6), data_in(5) => NPC1_IN(5), data_in(4) => 
                           NPC1_IN(4), data_in(3) => NPC1_IN(3), data_in(2) => 
                           NPC1_IN(2), data_in(1) => NPC1_IN(1), data_in(0) => 
                           NPC1_IN(0), data_out(31) => NPC1_OUT(31), 
                           data_out(30) => NPC1_OUT(30), data_out(29) => 
                           NPC1_OUT(29), data_out(28) => NPC1_OUT(28), 
                           data_out(27) => NPC1_OUT(27), data_out(26) => 
                           NPC1_OUT(26), data_out(25) => NPC1_OUT(25), 
                           data_out(24) => NPC1_OUT(24), data_out(23) => 
                           NPC1_OUT(23), data_out(22) => NPC1_OUT(22), 
                           data_out(21) => NPC1_OUT(21), data_out(20) => 
                           NPC1_OUT(20), data_out(19) => NPC1_OUT(19), 
                           data_out(18) => NPC1_OUT(18), data_out(17) => 
                           NPC1_OUT(17), data_out(16) => NPC1_OUT(16), 
                           data_out(15) => NPC1_OUT(15), data_out(14) => 
                           NPC1_OUT(14), data_out(13) => NPC1_OUT(13), 
                           data_out(12) => NPC1_OUT(12), data_out(11) => 
                           NPC1_OUT(11), data_out(10) => NPC1_OUT(10), 
                           data_out(9) => NPC1_OUT(9), data_out(8) => 
                           NPC1_OUT(8), data_out(7) => NPC1_OUT(7), data_out(6)
                           => NPC1_OUT(6), data_out(5) => NPC1_OUT(5), 
                           data_out(4) => NPC1_OUT(4), data_out(3) => 
                           NPC1_OUT(3), data_out(2) => NPC1_OUT(2), data_out(1)
                           => NPC1_OUT(1), data_out(0) => NPC1_OUT(0));
   IMM : gen_reg_N32_7 port map( clk => CLK, rst => RST, ld => DEC_OUTREG_EN, 
                           data_in(31) => SIGN_EXT_OUT_31_port, data_in(30) => 
                           SIGN_EXT_OUT_30_port, data_in(29) => 
                           SIGN_EXT_OUT_29_port, data_in(28) => 
                           SIGN_EXT_OUT_28_port, data_in(27) => 
                           SIGN_EXT_OUT_27_port, data_in(26) => 
                           SIGN_EXT_OUT_26_port, data_in(25) => 
                           SIGN_EXT_OUT_25_port, data_in(24) => 
                           SIGN_EXT_OUT_24_port, data_in(23) => 
                           SIGN_EXT_OUT_23_port, data_in(22) => 
                           SIGN_EXT_OUT_22_port, data_in(21) => 
                           SIGN_EXT_OUT_21_port, data_in(20) => 
                           SIGN_EXT_OUT_20_port, data_in(19) => 
                           SIGN_EXT_OUT_19_port, data_in(18) => 
                           SIGN_EXT_OUT_18_port, data_in(17) => 
                           SIGN_EXT_OUT_17_port, data_in(16) => 
                           SIGN_EXT_OUT_16_port, data_in(15) => 
                           SIGN_EXT_OUT_15_port, data_in(14) => 
                           SIGN_EXT_OUT_14_port, data_in(13) => 
                           SIGN_EXT_OUT_13_port, data_in(12) => 
                           SIGN_EXT_OUT_12_port, data_in(11) => 
                           SIGN_EXT_OUT_11_port, data_in(10) => 
                           SIGN_EXT_OUT_10_port, data_in(9) => 
                           SIGN_EXT_OUT_9_port, data_in(8) => 
                           SIGN_EXT_OUT_8_port, data_in(7) => 
                           SIGN_EXT_OUT_7_port, data_in(6) => 
                           SIGN_EXT_OUT_6_port, data_in(5) => 
                           SIGN_EXT_OUT_5_port, data_in(4) => 
                           SIGN_EXT_OUT_4_port, data_in(3) => 
                           SIGN_EXT_OUT_3_port, data_in(2) => 
                           SIGN_EXT_OUT_2_port, data_in(1) => 
                           SIGN_EXT_OUT_1_port, data_in(0) => 
                           SIGN_EXT_OUT_0_port, data_out(31) => REGIMM_OUT(31),
                           data_out(30) => REGIMM_OUT(30), data_out(29) => 
                           REGIMM_OUT(29), data_out(28) => REGIMM_OUT(28), 
                           data_out(27) => REGIMM_OUT(27), data_out(26) => 
                           REGIMM_OUT(26), data_out(25) => REGIMM_OUT(25), 
                           data_out(24) => REGIMM_OUT(24), data_out(23) => 
                           REGIMM_OUT(23), data_out(22) => REGIMM_OUT(22), 
                           data_out(21) => REGIMM_OUT(21), data_out(20) => 
                           REGIMM_OUT(20), data_out(19) => REGIMM_OUT(19), 
                           data_out(18) => REGIMM_OUT(18), data_out(17) => 
                           REGIMM_OUT(17), data_out(16) => REGIMM_OUT(16), 
                           data_out(15) => REGIMM_OUT(15), data_out(14) => 
                           REGIMM_OUT(14), data_out(13) => REGIMM_OUT(13), 
                           data_out(12) => REGIMM_OUT(12), data_out(11) => 
                           REGIMM_OUT(11), data_out(10) => REGIMM_OUT(10), 
                           data_out(9) => REGIMM_OUT(9), data_out(8) => 
                           REGIMM_OUT(8), data_out(7) => REGIMM_OUT(7), 
                           data_out(6) => REGIMM_OUT(6), data_out(5) => 
                           REGIMM_OUT(5), data_out(4) => REGIMM_OUT(4), 
                           data_out(3) => REGIMM_OUT(3), data_out(2) => 
                           REGIMM_OUT(2), data_out(1) => REGIMM_OUT(1), 
                           data_out(0) => REGIMM_OUT(0));
   WR_ADDR : gen_reg_N5_0 port map( clk => CLK, rst => RST, ld => DEC_OUTREG_EN
                           , data_in(4) => MUX_OUT_4_port, data_in(3) => 
                           MUX_OUT_3_port, data_in(2) => MUX_OUT_2_port, 
                           data_in(1) => MUX_OUT_1_port, data_in(0) => 
                           MUX_OUT_0_port, data_out(4) => WR_ADDR_OUT(4), 
                           data_out(3) => WR_ADDR_OUT(3), data_out(2) => 
                           WR_ADDR_OUT(2), data_out(1) => WR_ADDR_OUT(1), 
                           data_out(0) => WR_ADDR_OUT(0));
   RF : reg_file_Dbits32_Abits5 port map( CLK => CLK, RESET => RST, ENABLE => 
                           DEC_OUTREG_EN, RD1 => RD1_EN, RD2 => RD2_EN, WR => 
                           WR_EN, ADD_WR(4) => ADD_WR_4_port, ADD_WR(3) => 
                           ADD_WR_3_port, ADD_WR(2) => ADD_WR_2_port, ADD_WR(1)
                           => ADD_WR_1_port, ADD_WR(0) => ADD_WR_0_port, 
                           ADD_RD1(4) => I_CODE(25), ADD_RD1(3) => I_CODE(24), 
                           ADD_RD1(2) => I_CODE(23), ADD_RD1(1) => I_CODE(22), 
                           ADD_RD1(0) => I_CODE(21), ADD_RD2(4) => I_CODE(20), 
                           ADD_RD2(3) => I_CODE(19), ADD_RD2(2) => I_CODE(18), 
                           ADD_RD2(1) => I_CODE(17), ADD_RD2(0) => I_CODE(16), 
                           DATAIN(31) => DATA_IN(31), DATAIN(30) => DATA_IN(30)
                           , DATAIN(29) => DATA_IN(29), DATAIN(28) => 
                           DATA_IN(28), DATAIN(27) => DATA_IN(27), DATAIN(26) 
                           => DATA_IN(26), DATAIN(25) => DATA_IN(25), 
                           DATAIN(24) => DATA_IN(24), DATAIN(23) => DATA_IN(23)
                           , DATAIN(22) => DATA_IN(22), DATAIN(21) => 
                           DATA_IN(21), DATAIN(20) => DATA_IN(20), DATAIN(19) 
                           => DATA_IN(19), DATAIN(18) => DATA_IN(18), 
                           DATAIN(17) => DATA_IN(17), DATAIN(16) => DATA_IN(16)
                           , DATAIN(15) => DATA_IN(15), DATAIN(14) => 
                           DATA_IN(14), DATAIN(13) => DATA_IN(13), DATAIN(12) 
                           => DATA_IN(12), DATAIN(11) => DATA_IN(11), 
                           DATAIN(10) => DATA_IN(10), DATAIN(9) => DATA_IN(9), 
                           DATAIN(8) => DATA_IN(8), DATAIN(7) => DATA_IN(7), 
                           DATAIN(6) => DATA_IN(6), DATAIN(5) => DATA_IN(5), 
                           DATAIN(4) => DATA_IN(4), DATAIN(3) => DATA_IN(3), 
                           DATAIN(2) => DATA_IN(2), DATAIN(1) => DATA_IN(1), 
                           DATAIN(0) => DATA_IN(0), OUT1(31) => REGA_OUT(31), 
                           OUT1(30) => REGA_OUT(30), OUT1(29) => REGA_OUT(29), 
                           OUT1(28) => REGA_OUT(28), OUT1(27) => REGA_OUT(27), 
                           OUT1(26) => REGA_OUT(26), OUT1(25) => REGA_OUT(25), 
                           OUT1(24) => REGA_OUT(24), OUT1(23) => REGA_OUT(23), 
                           OUT1(22) => REGA_OUT(22), OUT1(21) => REGA_OUT(21), 
                           OUT1(20) => REGA_OUT(20), OUT1(19) => REGA_OUT(19), 
                           OUT1(18) => REGA_OUT(18), OUT1(17) => REGA_OUT(17), 
                           OUT1(16) => REGA_OUT(16), OUT1(15) => REGA_OUT(15), 
                           OUT1(14) => REGA_OUT(14), OUT1(13) => REGA_OUT(13), 
                           OUT1(12) => REGA_OUT(12), OUT1(11) => REGA_OUT(11), 
                           OUT1(10) => REGA_OUT(10), OUT1(9) => REGA_OUT(9), 
                           OUT1(8) => REGA_OUT(8), OUT1(7) => REGA_OUT(7), 
                           OUT1(6) => REGA_OUT(6), OUT1(5) => REGA_OUT(5), 
                           OUT1(4) => REGA_OUT(4), OUT1(3) => REGA_OUT(3), 
                           OUT1(2) => REGA_OUT(2), OUT1(1) => REGA_OUT(1), 
                           OUT1(0) => REGA_OUT(0), OUT2(31) => REGB_OUT(31), 
                           OUT2(30) => REGB_OUT(30), OUT2(29) => REGB_OUT(29), 
                           OUT2(28) => REGB_OUT(28), OUT2(27) => REGB_OUT(27), 
                           OUT2(26) => REGB_OUT(26), OUT2(25) => REGB_OUT(25), 
                           OUT2(24) => REGB_OUT(24), OUT2(23) => REGB_OUT(23), 
                           OUT2(22) => REGB_OUT(22), OUT2(21) => REGB_OUT(21), 
                           OUT2(20) => REGB_OUT(20), OUT2(19) => REGB_OUT(19), 
                           OUT2(18) => REGB_OUT(18), OUT2(17) => REGB_OUT(17), 
                           OUT2(16) => REGB_OUT(16), OUT2(15) => REGB_OUT(15), 
                           OUT2(14) => REGB_OUT(14), OUT2(13) => REGB_OUT(13), 
                           OUT2(12) => REGB_OUT(12), OUT2(11) => REGB_OUT(11), 
                           OUT2(10) => REGB_OUT(10), OUT2(9) => REGB_OUT(9), 
                           OUT2(8) => REGB_OUT(8), OUT2(7) => REGB_OUT(7), 
                           OUT2(6) => REGB_OUT(6), OUT2(5) => REGB_OUT(5), 
                           OUT2(4) => REGB_OUT(4), OUT2(3) => REGB_OUT(3), 
                           OUT2(2) => REGB_OUT(2), OUT2(1) => REGB_OUT(1), 
                           OUT2(0) => REGB_OUT(0));
   SING_EXT : sign_ext_N_IN026_N_IN116_N_OUT32 port map( ctrl_in => IS_I_TYPE, 
                           zero_padding => ZERO_PADDING2, data_in(25) => 
                           I_CODE(25), data_in(24) => I_CODE(24), data_in(23) 
                           => I_CODE(23), data_in(22) => I_CODE(22), 
                           data_in(21) => I_CODE(21), data_in(20) => I_CODE(20)
                           , data_in(19) => I_CODE(19), data_in(18) => 
                           I_CODE(18), data_in(17) => I_CODE(17), data_in(16) 
                           => I_CODE(16), data_in(15) => I_CODE(15), 
                           data_in(14) => I_CODE(14), data_in(13) => I_CODE(13)
                           , data_in(12) => I_CODE(12), data_in(11) => 
                           I_CODE(11), data_in(10) => I_CODE(10), data_in(9) =>
                           I_CODE(9), data_in(8) => I_CODE(8), data_in(7) => 
                           I_CODE(7), data_in(6) => I_CODE(6), data_in(5) => 
                           I_CODE(5), data_in(4) => I_CODE(4), data_in(3) => 
                           I_CODE(3), data_in(2) => I_CODE(2), data_in(1) => 
                           I_CODE(1), data_in(0) => I_CODE(0), data_ext(31) => 
                           SIGN_EXT_OUT_31_port, data_ext(30) => 
                           SIGN_EXT_OUT_30_port, data_ext(29) => 
                           SIGN_EXT_OUT_29_port, data_ext(28) => 
                           SIGN_EXT_OUT_28_port, data_ext(27) => 
                           SIGN_EXT_OUT_27_port, data_ext(26) => 
                           SIGN_EXT_OUT_26_port, data_ext(25) => 
                           SIGN_EXT_OUT_25_port, data_ext(24) => 
                           SIGN_EXT_OUT_24_port, data_ext(23) => 
                           SIGN_EXT_OUT_23_port, data_ext(22) => 
                           SIGN_EXT_OUT_22_port, data_ext(21) => 
                           SIGN_EXT_OUT_21_port, data_ext(20) => 
                           SIGN_EXT_OUT_20_port, data_ext(19) => 
                           SIGN_EXT_OUT_19_port, data_ext(18) => 
                           SIGN_EXT_OUT_18_port, data_ext(17) => 
                           SIGN_EXT_OUT_17_port, data_ext(16) => 
                           SIGN_EXT_OUT_16_port, data_ext(15) => 
                           SIGN_EXT_OUT_15_port, data_ext(14) => 
                           SIGN_EXT_OUT_14_port, data_ext(13) => 
                           SIGN_EXT_OUT_13_port, data_ext(12) => 
                           SIGN_EXT_OUT_12_port, data_ext(11) => 
                           SIGN_EXT_OUT_11_port, data_ext(10) => 
                           SIGN_EXT_OUT_10_port, data_ext(9) => 
                           SIGN_EXT_OUT_9_port, data_ext(8) => 
                           SIGN_EXT_OUT_8_port, data_ext(7) => 
                           SIGN_EXT_OUT_7_port, data_ext(6) => 
                           SIGN_EXT_OUT_6_port, data_ext(5) => 
                           SIGN_EXT_OUT_5_port, data_ext(4) => 
                           SIGN_EXT_OUT_4_port, data_ext(3) => 
                           SIGN_EXT_OUT_3_port, data_ext(2) => 
                           SIGN_EXT_OUT_2_port, data_ext(1) => 
                           SIGN_EXT_OUT_1_port, data_ext(0) => 
                           SIGN_EXT_OUT_0_port);
   MUX_WR_ADDR : gen_mux21_N5 port map( sel => IS_I_TYPE, x(4) => I_CODE(15), 
                           x(3) => I_CODE(14), x(2) => I_CODE(13), x(1) => 
                           I_CODE(12), x(0) => I_CODE(11), y(4) => I_CODE(20), 
                           y(3) => I_CODE(19), y(2) => I_CODE(18), y(1) => 
                           I_CODE(17), y(0) => I_CODE(16), m(4) => 
                           MUX_OUT_4_port, m(3) => MUX_OUT_3_port, m(2) => 
                           MUX_OUT_2_port, m(1) => MUX_OUT_1_port, m(0) => 
                           MUX_OUT_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity IF_STAGE_N_BITS_DATA32_N_BYTES_INST4 is

   port( CLK, RST, IF_LATCH_EN, PC_LATCH_EN : in std_logic;  PC_IN, IR_IN : in 
         std_logic_vector (31 downto 0);  PC_OUT, IR_OUT, NPC_OUT : out 
         std_logic_vector (31 downto 0));

end IF_STAGE_N_BITS_DATA32_N_BYTES_INST4;

architecture SYN_STRUCTURAL of IF_STAGE_N_BITS_DATA32_N_BYTES_INST4 is

   component pc_add_N32_OP24
      port( data_in : in std_logic_vector (31 downto 0);  data_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N32_9
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N32_10
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component gen_reg_N32_0
      port( clk, rst, ld : in std_logic;  data_in : in std_logic_vector (31 
            downto 0);  data_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal PC_OUT_31_port, PC_OUT_30_port, PC_OUT_29_port, PC_OUT_28_port, 
      PC_OUT_27_port, PC_OUT_26_port, PC_OUT_25_port, PC_OUT_24_port, 
      PC_OUT_23_port, PC_OUT_22_port, PC_OUT_21_port, PC_OUT_20_port, 
      PC_OUT_19_port, PC_OUT_18_port, PC_OUT_17_port, PC_OUT_16_port, 
      PC_OUT_15_port, PC_OUT_14_port, PC_OUT_13_port, PC_OUT_12_port, 
      PC_OUT_11_port, PC_OUT_10_port, PC_OUT_9_port, PC_OUT_8_port, 
      PC_OUT_7_port, PC_OUT_6_port, PC_OUT_5_port, PC_OUT_4_port, PC_OUT_3_port
      , PC_OUT_2_port, PC_OUT_1_port, PC_OUT_0_port, ADDER_OUT_31_port, 
      ADDER_OUT_30_port, ADDER_OUT_29_port, ADDER_OUT_28_port, 
      ADDER_OUT_27_port, ADDER_OUT_26_port, ADDER_OUT_25_port, 
      ADDER_OUT_24_port, ADDER_OUT_23_port, ADDER_OUT_22_port, 
      ADDER_OUT_21_port, ADDER_OUT_20_port, ADDER_OUT_19_port, 
      ADDER_OUT_18_port, ADDER_OUT_17_port, ADDER_OUT_16_port, 
      ADDER_OUT_15_port, ADDER_OUT_14_port, ADDER_OUT_13_port, 
      ADDER_OUT_12_port, ADDER_OUT_11_port, ADDER_OUT_10_port, ADDER_OUT_9_port
      , ADDER_OUT_8_port, ADDER_OUT_7_port, ADDER_OUT_6_port, ADDER_OUT_5_port,
      ADDER_OUT_4_port, ADDER_OUT_3_port, ADDER_OUT_2_port, ADDER_OUT_1_port, 
      ADDER_OUT_0_port : std_logic;

begin
   PC_OUT <= ( PC_OUT_31_port, PC_OUT_30_port, PC_OUT_29_port, PC_OUT_28_port, 
      PC_OUT_27_port, PC_OUT_26_port, PC_OUT_25_port, PC_OUT_24_port, 
      PC_OUT_23_port, PC_OUT_22_port, PC_OUT_21_port, PC_OUT_20_port, 
      PC_OUT_19_port, PC_OUT_18_port, PC_OUT_17_port, PC_OUT_16_port, 
      PC_OUT_15_port, PC_OUT_14_port, PC_OUT_13_port, PC_OUT_12_port, 
      PC_OUT_11_port, PC_OUT_10_port, PC_OUT_9_port, PC_OUT_8_port, 
      PC_OUT_7_port, PC_OUT_6_port, PC_OUT_5_port, PC_OUT_4_port, PC_OUT_3_port
      , PC_OUT_2_port, PC_OUT_1_port, PC_OUT_0_port );
   
   PC : gen_reg_N32_0 port map( clk => CLK, rst => RST, ld => PC_LATCH_EN, 
                           data_in(31) => PC_IN(31), data_in(30) => PC_IN(30), 
                           data_in(29) => PC_IN(29), data_in(28) => PC_IN(28), 
                           data_in(27) => PC_IN(27), data_in(26) => PC_IN(26), 
                           data_in(25) => PC_IN(25), data_in(24) => PC_IN(24), 
                           data_in(23) => PC_IN(23), data_in(22) => PC_IN(22), 
                           data_in(21) => PC_IN(21), data_in(20) => PC_IN(20), 
                           data_in(19) => PC_IN(19), data_in(18) => PC_IN(18), 
                           data_in(17) => PC_IN(17), data_in(16) => PC_IN(16), 
                           data_in(15) => PC_IN(15), data_in(14) => PC_IN(14), 
                           data_in(13) => PC_IN(13), data_in(12) => PC_IN(12), 
                           data_in(11) => PC_IN(11), data_in(10) => PC_IN(10), 
                           data_in(9) => PC_IN(9), data_in(8) => PC_IN(8), 
                           data_in(7) => PC_IN(7), data_in(6) => PC_IN(6), 
                           data_in(5) => PC_IN(5), data_in(4) => PC_IN(4), 
                           data_in(3) => PC_IN(3), data_in(2) => PC_IN(2), 
                           data_in(1) => PC_IN(1), data_in(0) => PC_IN(0), 
                           data_out(31) => PC_OUT_31_port, data_out(30) => 
                           PC_OUT_30_port, data_out(29) => PC_OUT_29_port, 
                           data_out(28) => PC_OUT_28_port, data_out(27) => 
                           PC_OUT_27_port, data_out(26) => PC_OUT_26_port, 
                           data_out(25) => PC_OUT_25_port, data_out(24) => 
                           PC_OUT_24_port, data_out(23) => PC_OUT_23_port, 
                           data_out(22) => PC_OUT_22_port, data_out(21) => 
                           PC_OUT_21_port, data_out(20) => PC_OUT_20_port, 
                           data_out(19) => PC_OUT_19_port, data_out(18) => 
                           PC_OUT_18_port, data_out(17) => PC_OUT_17_port, 
                           data_out(16) => PC_OUT_16_port, data_out(15) => 
                           PC_OUT_15_port, data_out(14) => PC_OUT_14_port, 
                           data_out(13) => PC_OUT_13_port, data_out(12) => 
                           PC_OUT_12_port, data_out(11) => PC_OUT_11_port, 
                           data_out(10) => PC_OUT_10_port, data_out(9) => 
                           PC_OUT_9_port, data_out(8) => PC_OUT_8_port, 
                           data_out(7) => PC_OUT_7_port, data_out(6) => 
                           PC_OUT_6_port, data_out(5) => PC_OUT_5_port, 
                           data_out(4) => PC_OUT_4_port, data_out(3) => 
                           PC_OUT_3_port, data_out(2) => PC_OUT_2_port, 
                           data_out(1) => PC_OUT_1_port, data_out(0) => 
                           PC_OUT_0_port);
   IR : gen_reg_N32_10 port map( clk => CLK, rst => RST, ld => IF_LATCH_EN, 
                           data_in(31) => IR_IN(31), data_in(30) => IR_IN(30), 
                           data_in(29) => IR_IN(29), data_in(28) => IR_IN(28), 
                           data_in(27) => IR_IN(27), data_in(26) => IR_IN(26), 
                           data_in(25) => IR_IN(25), data_in(24) => IR_IN(24), 
                           data_in(23) => IR_IN(23), data_in(22) => IR_IN(22), 
                           data_in(21) => IR_IN(21), data_in(20) => IR_IN(20), 
                           data_in(19) => IR_IN(19), data_in(18) => IR_IN(18), 
                           data_in(17) => IR_IN(17), data_in(16) => IR_IN(16), 
                           data_in(15) => IR_IN(15), data_in(14) => IR_IN(14), 
                           data_in(13) => IR_IN(13), data_in(12) => IR_IN(12), 
                           data_in(11) => IR_IN(11), data_in(10) => IR_IN(10), 
                           data_in(9) => IR_IN(9), data_in(8) => IR_IN(8), 
                           data_in(7) => IR_IN(7), data_in(6) => IR_IN(6), 
                           data_in(5) => IR_IN(5), data_in(4) => IR_IN(4), 
                           data_in(3) => IR_IN(3), data_in(2) => IR_IN(2), 
                           data_in(1) => IR_IN(1), data_in(0) => IR_IN(0), 
                           data_out(31) => IR_OUT(31), data_out(30) => 
                           IR_OUT(30), data_out(29) => IR_OUT(29), data_out(28)
                           => IR_OUT(28), data_out(27) => IR_OUT(27), 
                           data_out(26) => IR_OUT(26), data_out(25) => 
                           IR_OUT(25), data_out(24) => IR_OUT(24), data_out(23)
                           => IR_OUT(23), data_out(22) => IR_OUT(22), 
                           data_out(21) => IR_OUT(21), data_out(20) => 
                           IR_OUT(20), data_out(19) => IR_OUT(19), data_out(18)
                           => IR_OUT(18), data_out(17) => IR_OUT(17), 
                           data_out(16) => IR_OUT(16), data_out(15) => 
                           IR_OUT(15), data_out(14) => IR_OUT(14), data_out(13)
                           => IR_OUT(13), data_out(12) => IR_OUT(12), 
                           data_out(11) => IR_OUT(11), data_out(10) => 
                           IR_OUT(10), data_out(9) => IR_OUT(9), data_out(8) =>
                           IR_OUT(8), data_out(7) => IR_OUT(7), data_out(6) => 
                           IR_OUT(6), data_out(5) => IR_OUT(5), data_out(4) => 
                           IR_OUT(4), data_out(3) => IR_OUT(3), data_out(2) => 
                           IR_OUT(2), data_out(1) => IR_OUT(1), data_out(0) => 
                           IR_OUT(0));
   NPC : gen_reg_N32_9 port map( clk => CLK, rst => RST, ld => IF_LATCH_EN, 
                           data_in(31) => ADDER_OUT_31_port, data_in(30) => 
                           ADDER_OUT_30_port, data_in(29) => ADDER_OUT_29_port,
                           data_in(28) => ADDER_OUT_28_port, data_in(27) => 
                           ADDER_OUT_27_port, data_in(26) => ADDER_OUT_26_port,
                           data_in(25) => ADDER_OUT_25_port, data_in(24) => 
                           ADDER_OUT_24_port, data_in(23) => ADDER_OUT_23_port,
                           data_in(22) => ADDER_OUT_22_port, data_in(21) => 
                           ADDER_OUT_21_port, data_in(20) => ADDER_OUT_20_port,
                           data_in(19) => ADDER_OUT_19_port, data_in(18) => 
                           ADDER_OUT_18_port, data_in(17) => ADDER_OUT_17_port,
                           data_in(16) => ADDER_OUT_16_port, data_in(15) => 
                           ADDER_OUT_15_port, data_in(14) => ADDER_OUT_14_port,
                           data_in(13) => ADDER_OUT_13_port, data_in(12) => 
                           ADDER_OUT_12_port, data_in(11) => ADDER_OUT_11_port,
                           data_in(10) => ADDER_OUT_10_port, data_in(9) => 
                           ADDER_OUT_9_port, data_in(8) => ADDER_OUT_8_port, 
                           data_in(7) => ADDER_OUT_7_port, data_in(6) => 
                           ADDER_OUT_6_port, data_in(5) => ADDER_OUT_5_port, 
                           data_in(4) => ADDER_OUT_4_port, data_in(3) => 
                           ADDER_OUT_3_port, data_in(2) => ADDER_OUT_2_port, 
                           data_in(1) => ADDER_OUT_1_port, data_in(0) => 
                           ADDER_OUT_0_port, data_out(31) => NPC_OUT(31), 
                           data_out(30) => NPC_OUT(30), data_out(29) => 
                           NPC_OUT(29), data_out(28) => NPC_OUT(28), 
                           data_out(27) => NPC_OUT(27), data_out(26) => 
                           NPC_OUT(26), data_out(25) => NPC_OUT(25), 
                           data_out(24) => NPC_OUT(24), data_out(23) => 
                           NPC_OUT(23), data_out(22) => NPC_OUT(22), 
                           data_out(21) => NPC_OUT(21), data_out(20) => 
                           NPC_OUT(20), data_out(19) => NPC_OUT(19), 
                           data_out(18) => NPC_OUT(18), data_out(17) => 
                           NPC_OUT(17), data_out(16) => NPC_OUT(16), 
                           data_out(15) => NPC_OUT(15), data_out(14) => 
                           NPC_OUT(14), data_out(13) => NPC_OUT(13), 
                           data_out(12) => NPC_OUT(12), data_out(11) => 
                           NPC_OUT(11), data_out(10) => NPC_OUT(10), 
                           data_out(9) => NPC_OUT(9), data_out(8) => NPC_OUT(8)
                           , data_out(7) => NPC_OUT(7), data_out(6) => 
                           NPC_OUT(6), data_out(5) => NPC_OUT(5), data_out(4) 
                           => NPC_OUT(4), data_out(3) => NPC_OUT(3), 
                           data_out(2) => NPC_OUT(2), data_out(1) => NPC_OUT(1)
                           , data_out(0) => NPC_OUT(0));
   PC_ADDER : pc_add_N32_OP24 port map( data_in(31) => PC_OUT_31_port, 
                           data_in(30) => PC_OUT_30_port, data_in(29) => 
                           PC_OUT_29_port, data_in(28) => PC_OUT_28_port, 
                           data_in(27) => PC_OUT_27_port, data_in(26) => 
                           PC_OUT_26_port, data_in(25) => PC_OUT_25_port, 
                           data_in(24) => PC_OUT_24_port, data_in(23) => 
                           PC_OUT_23_port, data_in(22) => PC_OUT_22_port, 
                           data_in(21) => PC_OUT_21_port, data_in(20) => 
                           PC_OUT_20_port, data_in(19) => PC_OUT_19_port, 
                           data_in(18) => PC_OUT_18_port, data_in(17) => 
                           PC_OUT_17_port, data_in(16) => PC_OUT_16_port, 
                           data_in(15) => PC_OUT_15_port, data_in(14) => 
                           PC_OUT_14_port, data_in(13) => PC_OUT_13_port, 
                           data_in(12) => PC_OUT_12_port, data_in(11) => 
                           PC_OUT_11_port, data_in(10) => PC_OUT_10_port, 
                           data_in(9) => PC_OUT_9_port, data_in(8) => 
                           PC_OUT_8_port, data_in(7) => PC_OUT_7_port, 
                           data_in(6) => PC_OUT_6_port, data_in(5) => 
                           PC_OUT_5_port, data_in(4) => PC_OUT_4_port, 
                           data_in(3) => PC_OUT_3_port, data_in(2) => 
                           PC_OUT_2_port, data_in(1) => PC_OUT_1_port, 
                           data_in(0) => PC_OUT_0_port, data_out(31) => 
                           ADDER_OUT_31_port, data_out(30) => ADDER_OUT_30_port
                           , data_out(29) => ADDER_OUT_29_port, data_out(28) =>
                           ADDER_OUT_28_port, data_out(27) => ADDER_OUT_27_port
                           , data_out(26) => ADDER_OUT_26_port, data_out(25) =>
                           ADDER_OUT_25_port, data_out(24) => ADDER_OUT_24_port
                           , data_out(23) => ADDER_OUT_23_port, data_out(22) =>
                           ADDER_OUT_22_port, data_out(21) => ADDER_OUT_21_port
                           , data_out(20) => ADDER_OUT_20_port, data_out(19) =>
                           ADDER_OUT_19_port, data_out(18) => ADDER_OUT_18_port
                           , data_out(17) => ADDER_OUT_17_port, data_out(16) =>
                           ADDER_OUT_16_port, data_out(15) => ADDER_OUT_15_port
                           , data_out(14) => ADDER_OUT_14_port, data_out(13) =>
                           ADDER_OUT_13_port, data_out(12) => ADDER_OUT_12_port
                           , data_out(11) => ADDER_OUT_11_port, data_out(10) =>
                           ADDER_OUT_10_port, data_out(9) => ADDER_OUT_9_port, 
                           data_out(8) => ADDER_OUT_8_port, data_out(7) => 
                           ADDER_OUT_7_port, data_out(6) => ADDER_OUT_6_port, 
                           data_out(5) => ADDER_OUT_5_port, data_out(4) => 
                           ADDER_OUT_4_port, data_out(3) => ADDER_OUT_3_port, 
                           data_out(2) => ADDER_OUT_2_port, data_out(1) => 
                           ADDER_OUT_1_port, data_out(0) => ADDER_OUT_0_port);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE22 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, ZERO_PADDING2, 
         MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN : out std_logic;  
         ALU_OPCODE : out std_logic_vector (0 to 6);  FPU_OPCODE : out 
         std_logic_vector (0 to 4);  PC_LATCH_EN, MEM_OUTREG_EN, ZERO_PADDING4,
         MEM_OUT_SEL, DRAM_WE : out std_logic;  BYTE_LEN : out std_logic_vector
         (1 downto 0);  WB_MUX_SEL, JAL_MUX_SEL, WR_EN, WB_LATCH_EN : out 
         std_logic);

end CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE22;

architecture SYN_HARDWIRED of 
   CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFS_X1
      port( D, SI, SE, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, cw1_20_port, cw1_19_port, cw1_18_port, cw1_17_port, 
      cw1_16_port, cw1_15_port, cw1_14_port, cw1_13_port, cw1_12_port, 
      cw1_11_port, cw1_10_port, cw1_9_port, cw1_8_port, cw1_7_port, cw1_6_port,
      cw1_5_port, cw1_4_port, cw1_3_port, cw1_2_port, cw1_1_port, cw1_0_port, 
      cw2_15_port, cw2_14_port, cw2_13_port, cw2_12_port, cw2_11_port, 
      cw2_10_port, cw2_9_port, cw2_8_port, cw2_7_port, cw2_6_port, cw2_5_port, 
      cw2_4_port, cw2_3_port, cw2_2_port, cw2_1_port, cw2_0_port, cw3_10_port, 
      cw3_9_port, cw3_8_port, cw3_7_port, cw3_6_port, cw3_5_port, cw3_4_port, 
      cw3_3_port, cw3_2_port, cw3_1_port, cw3_0_port, cw4_3_port, cw4_2_port, 
      cw4_1_port, cw4_0_port, ALU_op1_6_port, ALU_op1_5_port, ALU_op1_4_port, 
      ALU_op1_3_port, ALU_op1_2_port, ALU_op1_1_port, ALU_op1_0_port, 
      ALU_op2_6_port, ALU_op2_5_port, ALU_op2_4_port, ALU_op2_3_port, 
      ALU_op2_2_port, ALU_op2_1_port, ALU_op2_0_port, FPU_op1_4_port, 
      FPU_op1_3_port, FPU_op1_2_port, FPU_op1_1_port, FPU_op1_0_port, 
      FPU_op2_4_port, FPU_op2_3_port, FPU_op2_2_port, FPU_op2_1_port, 
      FPU_op2_0_port, cw_18_port, cw_17_port, cw_16_port, cw_15_port, 
      cw_12_port, cw_11_port, cw_8_port, cw_5_port, cw_4_port, cw_3_port, 
      cw_2_port, ALU_op_5_port, n40, n48, n52, n59, n65, n84, n141, n142, n143,
      n144, n145, n300, n194, n54, n55, n56, n57, n58, n60, n61, n62, n63, n64,
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n134, n135, n136, n137, n138, n139, n140, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n195, n196, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n226, 
      n227, n228, n229, n230, n231, n232, n233, n237, n238, n236, n240, n255, 
      n256, n257, n258, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n284, n285, n286, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n301, n302, n303, n304, n306, n307, n308, 
      n309, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, 
      n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, 
      n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, 
      n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, 
      n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, 
      n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, 
      n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, 
      n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, 
      n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, 
      n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, 
      n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, 
      n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, 
      n_2205, n_2206, n_2207 : std_logic;

begin
   
   X_Logic1_port <= '1';
   n141 <= '0';
   n142 <= '1';
   n143 <= '1';
   n144 <= '1';
   n145 <= '0';
   U58 : AOI21_X1 port map( B1 => n270, B2 => n55, A => n194, ZN => n54);
   U59 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n84);
   U60 : AOI21_X1 port map( B1 => n58, B2 => n60, A => n260, ZN => n57);
   U61 : OAI21_X1 port map( B1 => n62, B2 => n261, A => IR_IN(27), ZN => n61);
   U62 : AOI21_X1 port map( B1 => n63, B2 => n64, A => IR_IN(28), ZN => n58);
   U63 : AOI22_X1 port map( A1 => n291, A2 => n66, B1 => n301, B2 => n67, ZN =>
                           n64);
   U64 : NOR2_X1 port map( A1 => n68, A2 => n307, ZN => n63);
   U65 : AOI22_X1 port map( A1 => IR_IN(31), A2 => n69, B1 => n70, B2 => n71, 
                           ZN => n56);
   U66 : OAI21_X1 port map( B1 => IR_IN(27), B2 => n72, A => n73, ZN => n69);
   U67 : NAND2_X1 port map( A1 => IR_IN(30), A2 => n273, ZN => n73);
   U68 : AOI22_X1 port map( A1 => n274, A2 => n271, B1 => n71, B2 => n279, ZN 
                           => n72);
   U69 : OR2_X1 port map( A1 => n74, A2 => n75, ZN => n65);
   U70 : OAI21_X1 port map( B1 => n276, B2 => n76, A => n77, ZN => n75);
   U71 : AOI22_X1 port map( A1 => n78, A2 => n275, B1 => n60, B2 => n70, ZN => 
                           n77);
   U72 : OAI21_X1 port map( B1 => n256, B2 => n277, A => n80, ZN => n74);
   U73 : AOI21_X1 port map( B1 => n81, B2 => n82, A => n83, ZN => n80);
   U74 : OAI21_X1 port map( B1 => n85, B2 => n261, A => n86, ZN => n59);
   U75 : AOI21_X1 port map( B1 => n87, B2 => n88, A => n262, ZN => n86);
   U76 : NAND2_X1 port map( A1 => IR_IN(28), A2 => n273, ZN => n88);
   U77 : AOI22_X1 port map( A1 => n90, A2 => n91, B1 => n92, B2 => IR_IN(29), 
                           ZN => n87);
   U78 : OAI21_X1 port map( B1 => n261, B2 => n281, A => IR_IN(28), ZN => n92);
   U79 : NOR3_X1 port map( A1 => n93, A2 => IR_IN(26), A3 => n94, ZN => n91);
   U80 : NOR3_X1 port map( A1 => n306, A2 => n95, A3 => n272, ZN => n90);
   U81 : AOI21_X1 port map( B1 => n96, B2 => n97, A => n285, ZN => n95);
   U82 : AOI22_X1 port map( A1 => n98, A2 => n99, B1 => IR_IN(30), B2 => n279, 
                           ZN => n85);
   U83 : NAND2_X1 port map( A1 => n79, A2 => IR_IN(26), ZN => n99);
   U84 : OAI21_X1 port map( B1 => n279, B2 => n100, A => IR_IN(29), ZN => n98);
   U85 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n270, ZN => n100);
   U86 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => n52);
   U87 : NOR3_X1 port map( A1 => n103, A2 => cw_8_port, A3 => n55, ZN => n102);
   U88 : NOR3_X1 port map( A1 => n277, A2 => n281, A3 => n256, ZN => n103);
   U89 : NOR3_X1 port map( A1 => n104, A2 => n105, A3 => n106, ZN => n101);
   U90 : NOR2_X1 port map( A1 => n107, A2 => n261, ZN => n106);
   U91 : AOI22_X1 port map( A1 => n79, A2 => n71, B1 => n108, B2 => n109, ZN =>
                           n107);
   U92 : NOR3_X1 port map( A1 => n110, A2 => IR_IN(31), A3 => IR_IN(28), ZN => 
                           n105);
   U93 : NOR2_X1 port map( A1 => n111, A2 => n265, ZN => n104);
   U94 : NOR3_X1 port map( A1 => n112, A2 => n293, A3 => n113, ZN => n111);
   U95 : OAI21_X1 port map( B1 => n115, B2 => n285, A => n116, ZN => n112);
   U96 : OR2_X1 port map( A1 => n117, A2 => n118, ZN => n48);
   U97 : OAI21_X1 port map( B1 => IR_IN(31), B2 => n282, A => n119, ZN => n118)
                           ;
   U98 : OAI21_X1 port map( B1 => n120, B2 => n121, A => IR_IN(31), ZN => n119)
                           ;
   U99 : OAI21_X1 port map( B1 => IR_IN(27), B2 => n122, A => n123, ZN => n121)
                           ;
   U100 : OAI21_X1 port map( B1 => n124, B2 => n62, A => IR_IN(27), ZN => n123)
                           ;
   U101 : OAI21_X1 port map( B1 => n125, B2 => n270, A => n126, ZN => n62);
   U102 : NAND2_X1 port map( A1 => n282, A2 => n273, ZN => n126);
   U103 : NOR2_X1 port map( A1 => n127, A2 => n271, ZN => n124);
   U104 : AOI22_X1 port map( A1 => n128, A2 => n271, B1 => n71, B2 => n280, ZN 
                           => n122);
   U105 : NOR2_X1 port map( A1 => IR_IN(29), A2 => n270, ZN => n120);
   U106 : OAI33_X1 port map( A1 => n264, A2 => n108, A3 => n281, B1 => n129, B2
                           => IR_IN(28), B3 => n130, ZN => n117);
   U107 : NOR3_X1 port map( A1 => n131, A2 => n132, A3 => n307, ZN => n130);
   U109 : AOI21_X1 port map( B1 => IR_IN(3), B2 => n137, A => IR_IN(26), ZN => 
                           n136);
   U110 : OAI21_X1 port map( B1 => n138, B2 => n139, A => n140, ZN => n134);
   U111 : AOI22_X1 port map( A1 => n146, A2 => n147, B1 => n298, B2 => n67, ZN 
                           => n140);
   U112 : NAND2_X1 port map( A1 => n148, A2 => n286, ZN => n131);
   U113 : AOI22_X1 port map( A1 => n150, A2 => n137, B1 => n302, B2 => n67, ZN 
                           => n148);
   U114 : OAI21_X1 port map( B1 => n151, B2 => n261, A => n152, ZN => n40);
   U115 : OAI21_X1 port map( B1 => n79, B2 => n269, A => n153, ZN => n152);
   U116 : OAI21_X1 port map( B1 => IR_IN(28), B2 => n129, A => n264, ZN => n153
                           );
   U117 : OAI21_X1 port map( B1 => n93, B2 => IR_IN(26), A => n270, ZN => n154)
                           ;
   U118 : NOR2_X1 port map( A1 => n155, A2 => n156, ZN => n93);
   U119 : OR2_X1 port map( A1 => n113, A2 => n82, ZN => n155);
   U120 : NAND2_X1 port map( A1 => n157, A2 => n116, ZN => n82);
   U121 : NOR4_X1 port map( A1 => n158, A2 => n135, A3 => n159, A4 => n132, ZN 
                           => n116);
   U122 : OAI21_X1 port map( B1 => n139, B2 => n96, A => n160, ZN => n132);
   U123 : AOI21_X1 port map( B1 => n161, B2 => n97, A => n139, ZN => n159);
   U124 : NOR2_X1 port map( A1 => n162, A2 => n139, ZN => n135);
   U125 : OR2_X1 port map( A1 => n163, A2 => n304, ZN => n162);
   U126 : NOR2_X1 port map( A1 => n291, A2 => n164, ZN => n157);
   U127 : NAND2_X1 port map( A1 => n150, A2 => n165, ZN => n139);
   U128 : AOI21_X1 port map( B1 => IR_IN(27), B2 => n277, A => n272, ZN => n151
                           );
   U129 : AOI21_X1 port map( B1 => IR_IN(26), B2 => IR_IN(28), A => n108, ZN =>
                           n128);
   U130 : AOI21_X1 port map( B1 => n267, B2 => n299, A => n166, ZN => n300);
   U131 : OAI21_X1 port map( B1 => n167, B2 => n168, A => n237, ZN => n166);
   U132 : NAND2_X1 port map( A1 => n169, A2 => n170, ZN => n237);
   U133 : NOR2_X1 port map( A1 => n297, A2 => n303, ZN => n167);
   U134 : NAND2_X1 port map( A1 => n171, A2 => n170, ZN => n168);
   U135 : NOR2_X1 port map( A1 => n172, A2 => n129, ZN => n170);
   U136 : NAND2_X1 port map( A1 => n125, A2 => n173, ZN => n172);
   U137 : NOR2_X1 port map( A1 => IR_IN(6), A2 => IR_IN(5), ZN => n171);
   U138 : NOR2_X1 port map( A1 => n255, A2 => n276, ZN => cw_8_port);
   U139 : NOR2_X1 port map( A1 => n281, A2 => n174, ZN => cw_5_port);
   U140 : OAI21_X1 port map( B1 => n282, B2 => n255, A => n174, ZN => cw_4_port
                           );
   U141 : NOR4_X1 port map( A1 => IR_IN(31), A2 => IR_IN(29), A3 => n280, A4 =>
                           n281, ZN => cw_2_port);
   U143 : NOR3_X1 port map( A1 => n76, A2 => n282, A3 => n281, ZN => n176);
   U144 : OAI21_X1 port map( B1 => n272, B2 => n179, A => n255, ZN => cw_3_port
                           );
   U145 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n125, ZN => n179);
   U146 : OR2_X1 port map( A1 => n266, A2 => n194, ZN => cw_18_port);
   U147 : NAND2_X1 port map( A1 => n180, A2 => n181, ZN => n194);
   U148 : AOI22_X1 port map( A1 => n182, A2 => n281, B1 => n263, B2 => n79, ZN 
                           => n180);
   U149 : OAI21_X1 port map( B1 => IR_IN(31), B2 => n274, A => n183, ZN => n182
                           );
   U150 : NAND2_X1 port map( A1 => n110, A2 => IR_IN(28), ZN => n183);
   U151 : OAI21_X1 port map( B1 => n76, B2 => n278, A => n184, ZN => cw_17_port
                           );
   U152 : NOR2_X1 port map( A1 => n238, A2 => n266, ZN => n184);
   U153 : NOR2_X1 port map( A1 => n186, A2 => n271, ZN => n238);
   U154 : OAI21_X1 port map( B1 => n187, B2 => n125, A => IR_IN(31), ZN => n186
                           );
   U155 : NOR2_X1 port map( A1 => IR_IN(28), A2 => IR_IN(27), ZN => n187);
   U156 : NAND2_X1 port map( A1 => n188, A2 => n189, ZN => cw_16_port);
   U157 : OAI21_X1 port map( B1 => n79, B2 => n127, A => n263, ZN => n189);
   U158 : NOR2_X1 port map( A1 => n281, A2 => n276, ZN => n79);
   U159 : AOI22_X1 port map( A1 => n190, A2 => n109, B1 => n191, B2 => n192, ZN
                           => n188);
   U160 : OAI21_X1 port map( B1 => n282, B2 => n281, A => n280, ZN => n192);
   U161 : NOR2_X1 port map( A1 => n193, A2 => n261, ZN => n190);
   U162 : NAND2_X1 port map( A1 => n195, A2 => n196, ZN => cw_15_port);
   U163 : AOI21_X1 port map( B1 => n263, B2 => IR_IN(27), A => n83, ZN => n196)
                           ;
   U164 : NOR2_X1 port map( A1 => n257, A2 => n178, ZN => n195);
   U165 : OAI21_X1 port map( B1 => n274, B2 => n76, A => n185, ZN => n178);
   U166 : OAI21_X1 port map( B1 => n156, B2 => n306, A => n81, ZN => n185);
   U167 : NOR2_X1 port map( A1 => n279, A2 => n129, ZN => n81);
   U169 : NAND2_X1 port map( A1 => n198, A2 => n199, ZN => n160);
   U170 : NOR3_X1 port map( A1 => n289, A2 => IR_IN(6), A3 => IR_IN(5), ZN => 
                           n199);
   U171 : NOR2_X1 port map( A1 => n296, A2 => n97, ZN => n198);
   U173 : NOR2_X1 port map( A1 => n201, A2 => n296, ZN => n150);
   U174 : NAND2_X1 port map( A1 => n295, A2 => IR_IN(5), ZN => n201);
   U175 : NOR2_X1 port map( A1 => n202, A2 => n292, ZN => n200);
   U176 : NOR2_X1 port map( A1 => n203, A2 => n202, ZN => n113);
   U178 : NOR2_X1 port map( A1 => n204, A2 => n302, ZN => n115);
   U179 : NAND2_X1 port map( A1 => n161, A2 => n205, ZN => n204);
   U180 : NOR2_X1 port map( A1 => n206, A2 => n97, ZN => n158);
   U181 : NAND2_X1 port map( A1 => n169, A2 => n67, ZN => n206);
   U182 : NAND2_X1 port map( A1 => n207, A2 => n208, ZN => n156);
   U183 : AOI21_X1 port map( B1 => n301, B2 => n290, A => n209, ZN => n208);
   U184 : NAND2_X1 port map( A1 => n210, A2 => n114, ZN => n209);
   U185 : NAND2_X1 port map( A1 => n211, A2 => n137, ZN => n114);
   U186 : NOR4_X1 port map( A1 => IR_IN(2), A2 => IR_IN(1), A3 => n294, A4 => 
                           n304, ZN => n137);
   U187 : NOR2_X1 port map( A1 => IR_IN(3), A2 => n212, ZN => n211);
   U188 : OAI21_X1 port map( B1 => n298, B2 => n147, A => n146, ZN => n210);
   U189 : NAND2_X1 port map( A1 => n213, A2 => IR_IN(0), ZN => n96);
   U190 : NOR2_X1 port map( A1 => IR_IN(1), A2 => n299, ZN => n213);
   U191 : NAND2_X1 port map( A1 => n147, A2 => IR_IN(2), ZN => n161);
   U192 : NOR2_X1 port map( A1 => IR_IN(1), A2 => IR_IN(0), ZN => n147);
   U193 : NOR2_X1 port map( A1 => n149, A2 => n68, ZN => n207);
   U194 : OAI21_X1 port map( B1 => n285, B2 => n138, A => n215, ZN => n68);
   U195 : NOR2_X1 port map( A1 => n94, A2 => n216, ZN => n215);
   U196 : NOR3_X1 port map( A1 => n304, A2 => n214, A3 => n163, ZN => n216);
   U197 : NOR2_X1 port map( A1 => n203, A2 => IR_IN(1), ZN => n94);
   U198 : OR2_X1 port map( A1 => n212, A2 => n292, ZN => n203);
   U199 : NOR2_X1 port map( A1 => n297, A2 => n294, ZN => n67);
   U200 : NAND2_X1 port map( A1 => n217, A2 => IR_IN(0), ZN => n138);
   U201 : NOR2_X1 port map( A1 => IR_IN(2), A2 => n303, ZN => n217);
   U202 : OAI21_X1 port map( B1 => n214, B2 => n97, A => n218, ZN => n149);
   U203 : NAND2_X1 port map( A1 => n146, A2 => n66, ZN => n218);
   U204 : NAND2_X1 port map( A1 => n97, A2 => n205, ZN => n66);
   U205 : NAND2_X1 port map( A1 => n219, A2 => IR_IN(1), ZN => n205);
   U206 : NOR2_X1 port map( A1 => IR_IN(2), A2 => IR_IN(0), ZN => n219);
   U207 : NOR2_X1 port map( A1 => n289, A2 => n212, ZN => n146);
   U208 : NAND2_X1 port map( A1 => n220, A2 => IR_IN(5), ZN => n212);
   U209 : NOR2_X1 port map( A1 => IR_IN(6), A2 => IR_IN(4), ZN => n220);
   U210 : OR2_X1 port map( A1 => n163, A2 => IR_IN(0), ZN => n97);
   U211 : NAND2_X1 port map( A1 => IR_IN(2), A2 => IR_IN(1), ZN => n163);
   U212 : NAND2_X1 port map( A1 => n165, A2 => n169, ZN => n214);
   U213 : NOR2_X1 port map( A1 => n221, A2 => IR_IN(4), ZN => n169);
   U214 : OR2_X1 port map( A1 => IR_IN(6), A2 => IR_IN(5), ZN => n221);
   U215 : NOR2_X1 port map( A1 => n294, A2 => IR_IN(3), ZN => n165);
   U216 : NOR4_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), A4 
                           => IR_IN(10), ZN => n173);
   U217 : NOR2_X1 port map( A1 => n222, A2 => n177, ZN => n181);
   U218 : OAI21_X1 port map( B1 => n193, B2 => n268, A => n223, ZN => n177);
   U219 : NOR2_X1 port map( A1 => n191, A2 => n224, ZN => n223);
   U220 : NOR3_X1 port map( A1 => n273, A2 => IR_IN(31), A3 => IR_IN(28), ZN =>
                           n224);
   U221 : AOI21_X1 port map( B1 => n281, B2 => IR_IN(28), A => n70, ZN => n193)
                           ;
   U222 : NAND2_X1 port map( A1 => n174, A2 => n309, ZN => n222);
   U224 : NAND2_X1 port map( A1 => n226, A2 => IR_IN(31), ZN => n174);
   U225 : NOR2_X1 port map( A1 => IR_IN(30), A2 => n280, ZN => n226);
   U226 : OAI21_X1 port map( B1 => n274, B2 => n129, A => n89, ZN => cw_12_port
                           );
   U227 : OAI21_X1 port map( B1 => n276, B2 => n129, A => n89, ZN => cw_11_port
                           );
   U228 : NAND2_X1 port map( A1 => n55, A2 => n273, ZN => n89);
   U229 : NOR2_X1 port map( A1 => n278, A2 => IR_IN(31), ZN => n55);
   U230 : NOR2_X1 port map( A1 => n281, A2 => IR_IN(28), ZN => n70);
   U231 : NAND2_X1 port map( A1 => n60, A2 => n281, ZN => n129);
   U232 : NAND2_X1 port map( A1 => n227, A2 => n228, ZN => ALU_op_5_port);
   U233 : NOR3_X1 port map( A1 => n83, A2 => n263, A3 => n191, ZN => n228);
   U234 : NOR2_X1 port map( A1 => n271, A2 => IR_IN(31), ZN => n191);
   U235 : NOR2_X1 port map( A1 => n273, A2 => IR_IN(30), ZN => n71);
   U236 : NAND2_X1 port map( A1 => n229, A2 => IR_IN(30), ZN => n76);
   U237 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(29), ZN => n229);
   U238 : NOR2_X1 port map( A1 => n256, A2 => IR_IN(27), ZN => n83);
   U239 : AOI21_X1 port map( B1 => n60, B2 => IR_IN(28), A => n231, ZN => n227)
                           ;
   U240 : OAI21_X1 port map( B1 => n232, B2 => n264, A => n233, ZN => n231);
   U241 : OAI21_X1 port map( B1 => n127, B2 => n125, A => n230, ZN => n233);
   U242 : NOR2_X1 port map( A1 => n272, A2 => n261, ZN => n230);
   U243 : NOR2_X1 port map( A1 => n276, A2 => IR_IN(26), ZN => n127);
   U244 : NOR2_X1 port map( A1 => n268, A2 => IR_IN(31), ZN => n78);
   U245 : NOR2_X1 port map( A1 => n270, A2 => n273, ZN => n109);
   U246 : NOR3_X1 port map( A1 => n281, A2 => n125, A3 => n108, ZN => n232);
   U247 : NOR2_X1 port map( A1 => IR_IN(28), A2 => IR_IN(26), ZN => n108);
   U248 : NOR2_X1 port map( A1 => n282, A2 => IR_IN(28), ZN => n125);
   U249 : NOR2_X1 port map( A1 => n272, A2 => IR_IN(31), ZN => n60);
   U250 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), ZN => n110);
   U9 : INV_X1 port map( A => n236, ZN => MUXA_SEL);
   U10 : INV_X1 port map( A => n240, ZN => MUXB_SEL);
   U11 : INV_X1 port map( A => n81, ZN => n265);
   U12 : INV_X1 port map( A => n185, ZN => n266);
   U13 : INV_X1 port map( A => n214, ZN => n290);
   U14 : INV_X1 port map( A => n146, ZN => n285);
   U15 : INV_X1 port map( A => n67, ZN => n292);
   U16 : INV_X1 port map( A => n139, ZN => n291);
   U17 : INV_X1 port map( A => n109, ZN => n268);
   U18 : INV_X1 port map( A => n230, ZN => n256);
   U19 : INV_X1 port map( A => n114, ZN => n293);
   U20 : INV_X1 port map( A => n149, ZN => n286);
   U21 : INV_X1 port map( A => n79, ZN => n275);
   U22 : INV_X1 port map( A => n125, ZN => n280);
   U23 : INV_X1 port map( A => n173, ZN => n294);
   U24 : INV_X1 port map( A => n71, ZN => n271);
   U25 : INV_X1 port map( A => n108, ZN => n279);
   U26 : INV_X1 port map( A => n127, ZN => n274);
   U27 : INV_X1 port map( A => n110, ZN => n272);
   U28 : INV_X1 port map( A => n76, ZN => n263);
   U29 : INV_X1 port map( A => n83, ZN => n255);
   U31 : INV_X1 port map( A => n160, ZN => n288);
   U33 : INV_X1 port map( A => n136, ZN => n284);
   U34 : INV_X1 port map( A => n168, ZN => n267);
   U36 : INV_X1 port map( A => n70, ZN => n278);
   U37 : INV_X1 port map( A => n128, ZN => n277);
   U38 : INV_X1 port map( A => n165, ZN => n289);
   U39 : INV_X1 port map( A => n78, ZN => n264);
   U40 : INV_X1 port map( A => n96, ZN => n298);
   U41 : INV_X1 port map( A => n161, ZN => n301);
   U42 : INV_X1 port map( A => n138, ZN => n302);
   U43 : INV_X1 port map( A => n54, ZN => n258);
   U44 : INV_X1 port map( A => IR_IN(6), ZN => n295);
   U45 : INV_X1 port map( A => IR_IN(27), ZN => n281);
   U47 : INV_X1 port map( A => IR_IN(29), ZN => n273);
   U48 : INV_X1 port map( A => IR_IN(31), ZN => n261);
   U49 : INV_X1 port map( A => n89, ZN => n262);
   U50 : INV_X1 port map( A => n154, ZN => n269);
   U51 : INV_X1 port map( A => IR_IN(30), ZN => n270);
   U52 : INV_X1 port map( A => IR_IN(26), ZN => n282);
   U53 : INV_X1 port map( A => IR_IN(28), ZN => n276);
   U54 : INV_X1 port map( A => n61, ZN => n260);
   U55 : INV_X1 port map( A => n181, ZN => n257);
   U56 : INV_X1 port map( A => IR_IN(0), ZN => n304);
   U57 : INV_X1 port map( A => IR_IN(3), ZN => n297);
   U251 : INV_X1 port map( A => IR_IN(4), ZN => n296);
   U252 : INV_X1 port map( A => IR_IN(2), ZN => n299);
   U253 : INV_X1 port map( A => IR_IN(1), ZN => n303);
   cw5_reg_0_inst : DFFR_X1 port map( D => cw4_0_port, CK => Clk, RN => Rst, Q 
                           => WB_LATCH_EN, QN => n_2098);
   cw3_reg_14_inst : DFFR_X1 port map( D => cw2_14_port, CK => Clk, RN => Rst, 
                           Q => n_2099, QN => n240);
   cw4_reg_10_inst : DFFR_X1 port map( D => cw3_10_port, CK => Clk, RN => Rst, 
                           Q => PC_LATCH_EN, QN => n_2100);
   cw3_reg_15_inst : DFFR_X1 port map( D => cw2_15_port, CK => Clk, RN => Rst, 
                           Q => n_2101, QN => n236);
   cw4_reg_7_inst : DFFR_X1 port map( D => cw3_7_port, CK => Clk, RN => Rst, Q 
                           => MEM_OUT_SEL, QN => n_2102);
   cw1_reg_21_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => Rst
                           , Q => IF_LATCH_EN, QN => n_2103);
   cw1_reg_20_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => Rst
                           , Q => cw1_20_port, QN => n_2104);
   cw1_reg_19_inst : DFFR_X1 port map( D => n194, CK => Clk, RN => Rst, Q => 
                           cw1_19_port, QN => n_2105);
   cw1_reg_18_inst : DFFR_X1 port map( D => cw_18_port, CK => Clk, RN => Rst, Q
                           => cw1_18_port, QN => n_2106);
   cw1_reg_17_inst : DFFR_X1 port map( D => cw_17_port, CK => Clk, RN => Rst, Q
                           => cw1_17_port, QN => n_2107);
   cw1_reg_16_inst : DFFR_X1 port map( D => cw_16_port, CK => Clk, RN => Rst, Q
                           => cw1_16_port, QN => n_2108);
   cw1_reg_15_inst : DFFR_X1 port map( D => cw_15_port, CK => Clk, RN => Rst, Q
                           => cw1_15_port, QN => n_2109);
   cw1_reg_14_inst : DFFR_X1 port map( D => n258, CK => Clk, RN => Rst, Q => 
                           cw1_14_port, QN => n_2110);
   cw1_reg_13_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => Rst
                           , Q => cw1_13_port, QN => n_2111);
   cw1_reg_12_inst : DFFR_X1 port map( D => cw_12_port, CK => Clk, RN => Rst, Q
                           => cw1_12_port, QN => n_2112);
   cw1_reg_11_inst : DFFR_X1 port map( D => cw_11_port, CK => Clk, RN => Rst, Q
                           => cw1_11_port, QN => n_2113);
   cw1_reg_10_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => Rst
                           , Q => cw1_10_port, QN => n_2114);
   cw1_reg_9_inst : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => Rst,
                           Q => cw1_9_port, QN => n_2115);
   cw1_reg_8_inst : DFFR_X1 port map( D => cw_8_port, CK => Clk, RN => Rst, Q 
                           => cw1_8_port, QN => n_2116);
   cw1_reg_7_inst : SDFFR_X1 port map( D => n145, SI => cw_5_port, SE => n273, 
                           CK => Clk, RN => Rst, Q => cw1_7_port, QN => n_2117)
                           ;
   cw1_reg_6_inst : DFFR_X1 port map( D => n238, CK => Clk, RN => Rst, Q => 
                           cw1_6_port, QN => n_2118);
   cw1_reg_5_inst : DFFR_X1 port map( D => cw_5_port, CK => Clk, RN => Rst, Q 
                           => cw1_5_port, QN => n_2119);
   cw1_reg_4_inst : DFFR_X1 port map( D => cw_4_port, CK => Clk, RN => Rst, Q 
                           => cw1_4_port, QN => n_2120);
   cw1_reg_3_inst : DFFR_X1 port map( D => cw_3_port, CK => Clk, RN => Rst, Q 
                           => cw1_3_port, QN => n_2121);
   cw1_reg_2_inst : DFFR_X1 port map( D => cw_2_port, CK => Clk, RN => Rst, Q 
                           => cw1_2_port, QN => n_2122);
   cw1_reg_1_inst : DFFR_X1 port map( D => n308, CK => Clk, RN => Rst, Q => 
                           cw1_1_port, QN => n_2123);
   cw1_reg_0_inst : DFFR_X1 port map( D => n308, CK => Clk, RN => Rst, Q => 
                           cw1_0_port, QN => n_2124);
   cw2_reg_20_inst : DFFR_X1 port map( D => cw1_20_port, CK => Clk, RN => Rst, 
                           Q => DEC_OUTREG_EN, QN => n_2125);
   cw2_reg_19_inst : DFFR_X1 port map( D => cw1_19_port, CK => Clk, RN => Rst, 
                           Q => IS_I_TYPE, QN => n_2126);
   cw2_reg_18_inst : DFFR_X1 port map( D => cw1_18_port, CK => Clk, RN => Rst, 
                           Q => RD1_EN, QN => n_2127);
   cw2_reg_17_inst : DFFR_X1 port map( D => cw1_17_port, CK => Clk, RN => Rst, 
                           Q => RD2_EN, QN => n_2128);
   cw2_reg_16_inst : DFFR_X1 port map( D => cw1_16_port, CK => Clk, RN => Rst, 
                           Q => ZERO_PADDING2, QN => n_2129);
   cw2_reg_15_inst : DFFR_X1 port map( D => cw1_15_port, CK => Clk, RN => Rst, 
                           Q => cw2_15_port, QN => n_2130);
   cw2_reg_14_inst : DFFR_X1 port map( D => cw1_14_port, CK => Clk, RN => Rst, 
                           Q => cw2_14_port, QN => n_2131);
   cw2_reg_13_inst : DFFR_X1 port map( D => cw1_13_port, CK => Clk, RN => Rst, 
                           Q => cw2_13_port, QN => n_2132);
   cw2_reg_12_inst : DFFR_X1 port map( D => cw1_12_port, CK => Clk, RN => Rst, 
                           Q => cw2_12_port, QN => n_2133);
   cw2_reg_11_inst : DFFR_X1 port map( D => cw1_11_port, CK => Clk, RN => Rst, 
                           Q => cw2_11_port, QN => n_2134);
   cw2_reg_10_inst : DFFR_X1 port map( D => cw1_10_port, CK => Clk, RN => Rst, 
                           Q => cw2_10_port, QN => n_2135);
   cw2_reg_9_inst : DFFR_X1 port map( D => cw1_9_port, CK => Clk, RN => Rst, Q 
                           => cw2_9_port, QN => n_2136);
   cw2_reg_8_inst : DFFR_X1 port map( D => cw1_8_port, CK => Clk, RN => Rst, Q 
                           => cw2_8_port, QN => n_2137);
   cw2_reg_7_inst : DFFR_X1 port map( D => cw1_7_port, CK => Clk, RN => Rst, Q 
                           => cw2_7_port, QN => n_2138);
   cw2_reg_6_inst : DFFR_X1 port map( D => cw1_6_port, CK => Clk, RN => Rst, Q 
                           => cw2_6_port, QN => n_2139);
   cw2_reg_5_inst : DFFR_X1 port map( D => cw1_5_port, CK => Clk, RN => Rst, Q 
                           => cw2_5_port, QN => n_2140);
   cw2_reg_4_inst : DFFR_X1 port map( D => cw1_4_port, CK => Clk, RN => Rst, Q 
                           => cw2_4_port, QN => n_2141);
   cw2_reg_3_inst : DFFR_X1 port map( D => cw1_3_port, CK => Clk, RN => Rst, Q 
                           => cw2_3_port, QN => n_2142);
   cw2_reg_2_inst : DFFR_X1 port map( D => cw1_2_port, CK => Clk, RN => Rst, Q 
                           => cw2_2_port, QN => n_2143);
   cw2_reg_1_inst : DFFR_X1 port map( D => cw1_1_port, CK => Clk, RN => Rst, Q 
                           => cw2_1_port, QN => n_2144);
   cw2_reg_0_inst : DFFR_X1 port map( D => cw1_0_port, CK => Clk, RN => Rst, Q 
                           => cw2_0_port, QN => n_2145);
   cw3_reg_13_inst : DFFR_X1 port map( D => cw2_13_port, CK => Clk, RN => Rst, 
                           Q => EXE_OUTREG_EN, QN => n_2146);
   cw3_reg_12_inst : DFFR_X1 port map( D => cw2_12_port, CK => Clk, RN => Rst, 
                           Q => EQ_COND, QN => n_2147);
   cw3_reg_11_inst : DFFR_X1 port map( D => cw2_11_port, CK => Clk, RN => Rst, 
                           Q => JUMP_EN, QN => n_2148);
   cw3_reg_10_inst : DFFR_X1 port map( D => cw2_10_port, CK => Clk, RN => Rst, 
                           Q => cw3_10_port, QN => n_2149);
   cw3_reg_9_inst : DFFR_X1 port map( D => cw2_9_port, CK => Clk, RN => Rst, Q 
                           => cw3_9_port, QN => n_2150);
   cw3_reg_8_inst : DFFR_X1 port map( D => cw2_8_port, CK => Clk, RN => Rst, Q 
                           => cw3_8_port, QN => n_2151);
   cw3_reg_7_inst : DFFR_X1 port map( D => cw2_7_port, CK => Clk, RN => Rst, Q 
                           => cw3_7_port, QN => n_2152);
   cw3_reg_6_inst : DFFR_X1 port map( D => cw2_6_port, CK => Clk, RN => Rst, Q 
                           => cw3_6_port, QN => n_2153);
   cw3_reg_5_inst : DFFR_X1 port map( D => cw2_5_port, CK => Clk, RN => Rst, Q 
                           => cw3_5_port, QN => n_2154);
   cw3_reg_4_inst : DFFR_X1 port map( D => cw2_4_port, CK => Clk, RN => Rst, Q 
                           => cw3_4_port, QN => n_2155);
   cw3_reg_3_inst : DFFR_X1 port map( D => cw2_3_port, CK => Clk, RN => Rst, Q 
                           => cw3_3_port, QN => n_2156);
   cw3_reg_2_inst : DFFR_X1 port map( D => cw2_2_port, CK => Clk, RN => Rst, Q 
                           => cw3_2_port, QN => n_2157);
   cw3_reg_1_inst : DFFR_X1 port map( D => cw2_1_port, CK => Clk, RN => Rst, Q 
                           => cw3_1_port, QN => n_2158);
   cw3_reg_0_inst : DFFR_X1 port map( D => cw2_0_port, CK => Clk, RN => Rst, Q 
                           => cw3_0_port, QN => n_2159);
   cw4_reg_9_inst : DFFR_X1 port map( D => cw3_9_port, CK => Clk, RN => Rst, Q 
                           => MEM_OUTREG_EN, QN => n_2160);
   cw4_reg_8_inst : DFFR_X1 port map( D => cw3_8_port, CK => Clk, RN => Rst, Q 
                           => ZERO_PADDING4, QN => n_2161);
   cw4_reg_6_inst : DFFR_X1 port map( D => cw3_6_port, CK => Clk, RN => Rst, Q 
                           => DRAM_WE, QN => n_2162);
   cw4_reg_5_inst : DFFR_X1 port map( D => cw3_5_port, CK => Clk, RN => Rst, Q 
                           => BYTE_LEN(1), QN => n_2163);
   cw4_reg_4_inst : DFFR_X1 port map( D => cw3_4_port, CK => Clk, RN => Rst, Q 
                           => BYTE_LEN(0), QN => n_2164);
   cw4_reg_3_inst : DFFR_X1 port map( D => cw3_3_port, CK => Clk, RN => Rst, Q 
                           => cw4_3_port, QN => n_2165);
   cw4_reg_2_inst : DFFR_X1 port map( D => cw3_2_port, CK => Clk, RN => Rst, Q 
                           => cw4_2_port, QN => n_2166);
   cw4_reg_1_inst : DFFR_X1 port map( D => cw3_1_port, CK => Clk, RN => Rst, Q 
                           => cw4_1_port, QN => n_2167);
   cw4_reg_0_inst : DFFR_X1 port map( D => cw3_0_port, CK => Clk, RN => Rst, Q 
                           => cw4_0_port, QN => n_2168);
   cw5_reg_3_inst : DFFR_X1 port map( D => cw4_3_port, CK => Clk, RN => Rst, Q 
                           => WB_MUX_SEL, QN => n_2169);
   cw5_reg_2_inst : DFFR_X1 port map( D => cw4_2_port, CK => Clk, RN => Rst, Q 
                           => JAL_MUX_SEL, QN => n_2170);
   cw5_reg_1_inst : DFFR_X1 port map( D => cw4_1_port, CK => Clk, RN => Rst, Q 
                           => WR_EN, QN => n_2171);
   ALU_op1_reg_6_inst : DFFS_X1 port map( D => n40, CK => Clk, SN => Rst, Q => 
                           ALU_op1_6_port, QN => n_2172);
   ALU_op1_reg_5_inst : DFFR_X1 port map( D => ALU_op_5_port, CK => Clk, RN => 
                           Rst, Q => ALU_op1_5_port, QN => n_2173);
   ALU_op1_reg_4_inst : DFFR_X1 port map( D => n65, CK => Clk, RN => Rst, Q => 
                           ALU_op1_4_port, QN => n_2174);
   ALU_op1_reg_3_inst : DFFS_X1 port map( D => n59, CK => Clk, SN => Rst, Q => 
                           ALU_op1_3_port, QN => n_2175);
   ALU_op1_reg_2_inst : DFFR_X1 port map( D => n52, CK => Clk, RN => Rst, Q => 
                           ALU_op1_2_port, QN => n_2176);
   ALU_op1_reg_1_inst : DFFS_X1 port map( D => n84, CK => Clk, SN => Rst, Q => 
                           ALU_op1_1_port, QN => n_2177);
   ALU_op1_reg_0_inst : DFFS_X1 port map( D => n48, CK => Clk, SN => Rst, Q => 
                           ALU_op1_0_port, QN => n_2178);
   ALU_op2_reg_5_inst : DFFR_X1 port map( D => ALU_op1_5_port, CK => Clk, RN =>
                           Rst, Q => ALU_op2_5_port, QN => n_2179);
   ALU_op2_reg_4_inst : DFFR_X1 port map( D => ALU_op1_4_port, CK => Clk, RN =>
                           Rst, Q => ALU_op2_4_port, QN => n_2180);
   ALU_op2_reg_2_inst : DFFR_X1 port map( D => ALU_op1_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_op2_2_port, QN => n_2181);
   ALU_op3_reg_5_inst : DFFR_X1 port map( D => ALU_op2_5_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPCODE(1), QN => n_2182);
   ALU_op3_reg_4_inst : DFFR_X1 port map( D => ALU_op2_4_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPCODE(2), QN => n_2183);
   ALU_op3_reg_2_inst : DFFR_X1 port map( D => ALU_op2_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPCODE(4), QN => n_2184);
   FPU_op1_reg_4_inst : DFFS_X1 port map( D => n237, CK => Clk, SN => Rst, Q =>
                           FPU_op1_4_port, QN => n_2185);
   FPU_op1_reg_3_inst : SDFFS_X1 port map( D => n144, SI => IR_IN(3), SE => 
                           n267, CK => Clk, SN => Rst, Q => FPU_op1_3_port, QN 
                           => n_2186);
   FPU_op1_reg_2_inst : SDFFS_X1 port map( D => n143, SI => IR_IN(2), SE => 
                           n267, CK => Clk, SN => Rst, Q => FPU_op1_2_port, QN 
                           => n_2187);
   FPU_op1_reg_1_inst : SDFFS_X1 port map( D => n142, SI => IR_IN(1), SE => 
                           n267, CK => Clk, SN => Rst, Q => FPU_op1_1_port, QN 
                           => n_2188);
   FPU_op1_reg_0_inst : SDFFR_X1 port map( D => IR_IN(0), SI => n141, SE => 
                           n300, CK => Clk, RN => Rst, Q => FPU_op1_0_port, QN 
                           => n_2189);
   FPU_op2_reg_0_inst : DFFR_X1 port map( D => FPU_op1_0_port, CK => Clk, RN =>
                           Rst, Q => FPU_op2_0_port, QN => n_2190);
   FPU_op3_reg_0_inst : DFFR_X1 port map( D => FPU_op2_0_port, CK => Clk, RN =>
                           Rst, Q => FPU_OPCODE(4), QN => n_2191);
   FPU_op2_reg_3_inst : DFFS_X1 port map( D => FPU_op1_3_port, CK => Clk, SN =>
                           Rst, Q => FPU_op2_3_port, QN => n_2192);
   FPU_op2_reg_2_inst : DFFS_X1 port map( D => FPU_op1_2_port, CK => Clk, SN =>
                           Rst, Q => FPU_op2_2_port, QN => n_2193);
   FPU_op2_reg_1_inst : DFFS_X1 port map( D => FPU_op1_1_port, CK => Clk, SN =>
                           Rst, Q => FPU_op2_1_port, QN => n_2194);
   FPU_op2_reg_4_inst : DFFS_X1 port map( D => FPU_op1_4_port, CK => Clk, SN =>
                           Rst, Q => FPU_op2_4_port, QN => n_2195);
   ALU_op3_reg_3_inst : DFFS_X1 port map( D => ALU_op2_3_port, CK => Clk, SN =>
                           Rst, Q => ALU_OPCODE(3), QN => n_2196);
   ALU_op2_reg_3_inst : DFFS_X1 port map( D => ALU_op1_3_port, CK => Clk, SN =>
                           Rst, Q => ALU_op2_3_port, QN => n_2197);
   FPU_op3_reg_4_inst : DFFS_X1 port map( D => FPU_op2_4_port, CK => Clk, SN =>
                           Rst, Q => FPU_OPCODE(0), QN => n_2198);
   FPU_op3_reg_3_inst : DFFS_X1 port map( D => FPU_op2_3_port, CK => Clk, SN =>
                           Rst, Q => FPU_OPCODE(1), QN => n_2199);
   FPU_op3_reg_2_inst : DFFS_X1 port map( D => FPU_op2_2_port, CK => Clk, SN =>
                           Rst, Q => FPU_OPCODE(2), QN => n_2200);
   FPU_op3_reg_1_inst : DFFS_X1 port map( D => FPU_op2_1_port, CK => Clk, SN =>
                           Rst, Q => FPU_OPCODE(3), QN => n_2201);
   ALU_op2_reg_6_inst : DFFS_X1 port map( D => ALU_op1_6_port, CK => Clk, SN =>
                           Rst, Q => ALU_op2_6_port, QN => n_2202);
   ALU_op2_reg_1_inst : DFFS_X1 port map( D => ALU_op1_1_port, CK => Clk, SN =>
                           Rst, Q => ALU_op2_1_port, QN => n_2203);
   ALU_op2_reg_0_inst : DFFS_X1 port map( D => ALU_op1_0_port, CK => Clk, SN =>
                           Rst, Q => ALU_op2_0_port, QN => n_2204);
   ALU_op3_reg_6_inst : DFFS_X1 port map( D => ALU_op2_6_port, CK => Clk, SN =>
                           Rst, Q => ALU_OPCODE(0), QN => n_2205);
   ALU_op3_reg_0_inst : DFFS_X1 port map( D => ALU_op2_0_port, CK => Clk, SN =>
                           Rst, Q => ALU_OPCODE(6), QN => n_2206);
   ALU_op3_reg_1_inst : DFFS_X1 port map( D => ALU_op2_1_port, CK => Clk, SN =>
                           Rst, Q => ALU_OPCODE(5), QN => n_2207);
   U8 : OR4_X1 port map( A1 => n158, A2 => n113, A3 => n164, A4 => n288, ZN => 
                           n306);
   U30 : OR4_X1 port map( A1 => n134, A2 => n284, A3 => n135, A4 => n93, ZN => 
                           n307);
   U32 : OR4_X1 port map( A1 => cw_3_port, A2 => n176, A3 => n177, A4 => n178, 
                           ZN => n308);
   U35 : OR4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(28), A3 => IR_IN(27), A4
                           => n261, ZN => n309);
   U46 : AND2_X1 port map( A1 => n115, A2 => n96, ZN => n202);
   U108 : AND2_X1 port map( A1 => n200, A2 => n150, ZN => n164);

end SYN_HARDWIRED;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 is

   port( CLK, RST, IF_LATCH_EN, PC_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, 
         RD2_EN, WR_EN, ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, 
         EQ_COND, JUMP_EN : in std_logic;  ALU_OPCODE : in std_logic_vector (0 
         to 6);  MEM_OUTREG_EN, ZERO_PADDING4, MEM_OUT_SEL : in std_logic;  
         BYTE_LEN_IN : in std_logic_vector (1 downto 0);  DRAM_WE : in 
         std_logic;  DRAM_WE_OUT : out std_logic;  BYTE_LEN_OUT : out 
         std_logic_vector (1 downto 0);  WB_LATCH_EN, JAL_MUX_SEL, WB_MUX_SEL :
         in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  PC_OUT : 
         out std_logic_vector (31 downto 0);  MEM_DATA_OUT_INT : in 
         std_logic_vector (31 downto 0);  MEM_ADDR_OUT, MEM_DATA_IN_PRIME : out
         std_logic_vector (31 downto 0));

end DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16;

architecture SYN_PIPELINED of 
   DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 is

   component WB_STAGE_N_BITS_DATA32_RF_ADDR5
      port( CLK, RST, WB_LATCH_EN, JAL_MUX_SEL, WB_MUX_SEL : in std_logic;  
            IR_IN : in std_logic_vector (4 downto 0);  MUX_IN2, MUX_IN1, 
            MUX_IN0 : in std_logic_vector (31 downto 0);  WRT_OUT : out 
            std_logic_vector (31 downto 0);  IR_OUT : out std_logic_vector (4 
            downto 0));
   end component;
   
   component MEM_STAGE_N_BITS_DATA32_RF_ADDR5
      port( CLK, RST, MEM_OUTREG_EN, ZERO_PADDING4, MEM_OUT_SEL : in std_logic;
            BYTE_LEN_IN : in std_logic_vector (1 downto 0);  DRAM_WE : in 
            std_logic;  DRAM_WE_OUT : out std_logic;  BYTE_LEN_OUT : out 
            std_logic_vector (1 downto 0);  BRA_IN : in std_logic;  
            JUMP_MUX_IN_0, ALU_OUTPUT_IN, MEM_DATA_IN, MEM_DATA_OUT_INT, NPC_IN
            : in std_logic_vector (31 downto 0);  IR_IN : in std_logic_vector 
            (4 downto 0);  IR_OUT : out std_logic_vector (4 downto 0);  NPC_OUT
            , MEM_ADDR_OUT, MEM_DATA_IN_PRIME, ALU_OUTPUT_OUT, MEM_DATA_OUT, 
            ADDR_MUX_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component EXE_STAGE_N_BITS_DATA32_RF_ADDR5
      port( CLK, RST, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN : in 
            std_logic;  ALU_OPCODE : in std_logic_vector (0 to 6);  NPC2_IN, 
            NPC1_MUXA_IN, REGA_MUXA_IN, REGB_MUXB_IN, IMM_MUXB_IN, PAD_IN : in 
            std_logic_vector (31 downto 0);  IR2_IN : in std_logic_vector (4 
            downto 0);  NPC2_OUT : out std_logic_vector (31 downto 0);  
            ZERO_OP_OUT : out std_logic;  ALU_OUT, PAD_OUT : out 
            std_logic_vector (31 downto 0);  IR2_OUT : out std_logic_vector (4 
            downto 0);  N_FLAG, Z_FLAG, C_FLAG, V_FLAG : out std_logic);
   end component;
   
   component 
      ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16
      port( CLK, RST, JAL_MUX_SEL, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, 
            WR_EN, ZERO_PADDING2 : in std_logic;  I_CODE, NPC1_IN, DATA_IN : in
            std_logic_vector (31 downto 0);  WR_ADDR_IN : in std_logic_vector 
            (4 downto 0);  REGA_OUT, REGB_OUT, REGIMM_OUT : out 
            std_logic_vector (31 downto 0);  WR_ADDR_OUT : out std_logic_vector
            (4 downto 0);  NPC1_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component IF_STAGE_N_BITS_DATA32_N_BYTES_INST4
      port( CLK, RST, IF_LATCH_EN, PC_LATCH_EN : in std_logic;  PC_IN, IR_IN : 
            in std_logic_vector (31 downto 0);  PC_OUT, IR_OUT, NPC_OUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal PC_MEM2IF_31_port, PC_MEM2IF_30_port, PC_MEM2IF_29_port, 
      PC_MEM2IF_28_port, PC_MEM2IF_27_port, PC_MEM2IF_26_port, 
      PC_MEM2IF_25_port, PC_MEM2IF_24_port, PC_MEM2IF_23_port, 
      PC_MEM2IF_22_port, PC_MEM2IF_21_port, PC_MEM2IF_20_port, 
      PC_MEM2IF_19_port, PC_MEM2IF_18_port, PC_MEM2IF_17_port, 
      PC_MEM2IF_16_port, PC_MEM2IF_15_port, PC_MEM2IF_14_port, 
      PC_MEM2IF_13_port, PC_MEM2IF_12_port, PC_MEM2IF_11_port, 
      PC_MEM2IF_10_port, PC_MEM2IF_9_port, PC_MEM2IF_8_port, PC_MEM2IF_7_port, 
      PC_MEM2IF_6_port, PC_MEM2IF_5_port, PC_MEM2IF_4_port, PC_MEM2IF_3_port, 
      PC_MEM2IF_2_port, PC_MEM2IF_1_port, PC_MEM2IF_0_port, IR_IF2ID_31_port, 
      IR_IF2ID_30_port, IR_IF2ID_29_port, IR_IF2ID_28_port, IR_IF2ID_27_port, 
      IR_IF2ID_26_port, IR_IF2ID_25_port, IR_IF2ID_24_port, IR_IF2ID_23_port, 
      IR_IF2ID_22_port, IR_IF2ID_21_port, IR_IF2ID_20_port, IR_IF2ID_19_port, 
      IR_IF2ID_18_port, IR_IF2ID_17_port, IR_IF2ID_16_port, IR_IF2ID_15_port, 
      IR_IF2ID_14_port, IR_IF2ID_13_port, IR_IF2ID_12_port, IR_IF2ID_11_port, 
      IR_IF2ID_10_port, IR_IF2ID_9_port, IR_IF2ID_8_port, IR_IF2ID_7_port, 
      IR_IF2ID_6_port, IR_IF2ID_5_port, IR_IF2ID_4_port, IR_IF2ID_3_port, 
      IR_IF2ID_2_port, IR_IF2ID_1_port, IR_IF2ID_0_port, NPC_IF2ID_MEM_31_port,
      NPC_IF2ID_MEM_30_port, NPC_IF2ID_MEM_29_port, NPC_IF2ID_MEM_28_port, 
      NPC_IF2ID_MEM_27_port, NPC_IF2ID_MEM_26_port, NPC_IF2ID_MEM_25_port, 
      NPC_IF2ID_MEM_24_port, NPC_IF2ID_MEM_23_port, NPC_IF2ID_MEM_22_port, 
      NPC_IF2ID_MEM_21_port, NPC_IF2ID_MEM_20_port, NPC_IF2ID_MEM_19_port, 
      NPC_IF2ID_MEM_18_port, NPC_IF2ID_MEM_17_port, NPC_IF2ID_MEM_16_port, 
      NPC_IF2ID_MEM_15_port, NPC_IF2ID_MEM_14_port, NPC_IF2ID_MEM_13_port, 
      NPC_IF2ID_MEM_12_port, NPC_IF2ID_MEM_11_port, NPC_IF2ID_MEM_10_port, 
      NPC_IF2ID_MEM_9_port, NPC_IF2ID_MEM_8_port, NPC_IF2ID_MEM_7_port, 
      NPC_IF2ID_MEM_6_port, NPC_IF2ID_MEM_5_port, NPC_IF2ID_MEM_4_port, 
      NPC_IF2ID_MEM_3_port, NPC_IF2ID_MEM_2_port, NPC_IF2ID_MEM_1_port, 
      NPC_IF2ID_MEM_0_port, WRT_WB2ID_31_port, WRT_WB2ID_30_port, 
      WRT_WB2ID_29_port, WRT_WB2ID_28_port, WRT_WB2ID_27_port, 
      WRT_WB2ID_26_port, WRT_WB2ID_25_port, WRT_WB2ID_24_port, 
      WRT_WB2ID_23_port, WRT_WB2ID_22_port, WRT_WB2ID_21_port, 
      WRT_WB2ID_20_port, WRT_WB2ID_19_port, WRT_WB2ID_18_port, 
      WRT_WB2ID_17_port, WRT_WB2ID_16_port, WRT_WB2ID_15_port, 
      WRT_WB2ID_14_port, WRT_WB2ID_13_port, WRT_WB2ID_12_port, 
      WRT_WB2ID_11_port, WRT_WB2ID_10_port, WRT_WB2ID_9_port, WRT_WB2ID_8_port,
      WRT_WB2ID_7_port, WRT_WB2ID_6_port, WRT_WB2ID_5_port, WRT_WB2ID_4_port, 
      WRT_WB2ID_3_port, WRT_WB2ID_2_port, WRT_WB2ID_1_port, WRT_WB2ID_0_port, 
      IR_WB2ID_4_port, IR_WB2ID_3_port, IR_WB2ID_2_port, IR_WB2ID_1_port, 
      IR_WB2ID_0_port, A_ID2EXE_31_port, A_ID2EXE_30_port, A_ID2EXE_29_port, 
      A_ID2EXE_28_port, A_ID2EXE_27_port, A_ID2EXE_26_port, A_ID2EXE_25_port, 
      A_ID2EXE_24_port, A_ID2EXE_23_port, A_ID2EXE_22_port, A_ID2EXE_21_port, 
      A_ID2EXE_20_port, A_ID2EXE_19_port, A_ID2EXE_18_port, A_ID2EXE_17_port, 
      A_ID2EXE_16_port, A_ID2EXE_15_port, A_ID2EXE_14_port, A_ID2EXE_13_port, 
      A_ID2EXE_12_port, A_ID2EXE_11_port, A_ID2EXE_10_port, A_ID2EXE_9_port, 
      A_ID2EXE_8_port, A_ID2EXE_7_port, A_ID2EXE_6_port, A_ID2EXE_5_port, 
      A_ID2EXE_4_port, A_ID2EXE_3_port, A_ID2EXE_2_port, A_ID2EXE_1_port, 
      A_ID2EXE_0_port, B_ID2EXE_31_port, B_ID2EXE_30_port, B_ID2EXE_29_port, 
      B_ID2EXE_28_port, B_ID2EXE_27_port, B_ID2EXE_26_port, B_ID2EXE_25_port, 
      B_ID2EXE_24_port, B_ID2EXE_23_port, B_ID2EXE_22_port, B_ID2EXE_21_port, 
      B_ID2EXE_20_port, B_ID2EXE_19_port, B_ID2EXE_18_port, B_ID2EXE_17_port, 
      B_ID2EXE_16_port, B_ID2EXE_15_port, B_ID2EXE_14_port, B_ID2EXE_13_port, 
      B_ID2EXE_12_port, B_ID2EXE_11_port, B_ID2EXE_10_port, B_ID2EXE_9_port, 
      B_ID2EXE_8_port, B_ID2EXE_7_port, B_ID2EXE_6_port, B_ID2EXE_5_port, 
      B_ID2EXE_4_port, B_ID2EXE_3_port, B_ID2EXE_2_port, B_ID2EXE_1_port, 
      B_ID2EXE_0_port, IMM_ID2EXE_31_port, IMM_ID2EXE_30_port, 
      IMM_ID2EXE_29_port, IMM_ID2EXE_28_port, IMM_ID2EXE_27_port, 
      IMM_ID2EXE_26_port, IMM_ID2EXE_25_port, IMM_ID2EXE_24_port, 
      IMM_ID2EXE_23_port, IMM_ID2EXE_22_port, IMM_ID2EXE_21_port, 
      IMM_ID2EXE_20_port, IMM_ID2EXE_19_port, IMM_ID2EXE_18_port, 
      IMM_ID2EXE_17_port, IMM_ID2EXE_16_port, IMM_ID2EXE_15_port, 
      IMM_ID2EXE_14_port, IMM_ID2EXE_13_port, IMM_ID2EXE_12_port, 
      IMM_ID2EXE_11_port, IMM_ID2EXE_10_port, IMM_ID2EXE_9_port, 
      IMM_ID2EXE_8_port, IMM_ID2EXE_7_port, IMM_ID2EXE_6_port, 
      IMM_ID2EXE_5_port, IMM_ID2EXE_4_port, IMM_ID2EXE_3_port, 
      IMM_ID2EXE_2_port, IMM_ID2EXE_1_port, IMM_ID2EXE_0_port, IR_ID2EXE_4_port
      , IR_ID2EXE_3_port, IR_ID2EXE_2_port, IR_ID2EXE_1_port, IR_ID2EXE_0_port,
      NPC_ID2EXE_31_port, NPC_ID2EXE_30_port, NPC_ID2EXE_29_port, 
      NPC_ID2EXE_28_port, NPC_ID2EXE_27_port, NPC_ID2EXE_26_port, 
      NPC_ID2EXE_25_port, NPC_ID2EXE_24_port, NPC_ID2EXE_23_port, 
      NPC_ID2EXE_22_port, NPC_ID2EXE_21_port, NPC_ID2EXE_20_port, 
      NPC_ID2EXE_19_port, NPC_ID2EXE_18_port, NPC_ID2EXE_17_port, 
      NPC_ID2EXE_16_port, NPC_ID2EXE_15_port, NPC_ID2EXE_14_port, 
      NPC_ID2EXE_13_port, NPC_ID2EXE_12_port, NPC_ID2EXE_11_port, 
      NPC_ID2EXE_10_port, NPC_ID2EXE_9_port, NPC_ID2EXE_8_port, 
      NPC_ID2EXE_7_port, NPC_ID2EXE_6_port, NPC_ID2EXE_5_port, 
      NPC_ID2EXE_4_port, NPC_ID2EXE_3_port, NPC_ID2EXE_2_port, 
      NPC_ID2EXE_1_port, NPC_ID2EXE_0_port, NPC_EXE2MEM_31_port, 
      NPC_EXE2MEM_30_port, NPC_EXE2MEM_29_port, NPC_EXE2MEM_28_port, 
      NPC_EXE2MEM_27_port, NPC_EXE2MEM_26_port, NPC_EXE2MEM_25_port, 
      NPC_EXE2MEM_24_port, NPC_EXE2MEM_23_port, NPC_EXE2MEM_22_port, 
      NPC_EXE2MEM_21_port, NPC_EXE2MEM_20_port, NPC_EXE2MEM_19_port, 
      NPC_EXE2MEM_18_port, NPC_EXE2MEM_17_port, NPC_EXE2MEM_16_port, 
      NPC_EXE2MEM_15_port, NPC_EXE2MEM_14_port, NPC_EXE2MEM_13_port, 
      NPC_EXE2MEM_12_port, NPC_EXE2MEM_11_port, NPC_EXE2MEM_10_port, 
      NPC_EXE2MEM_9_port, NPC_EXE2MEM_8_port, NPC_EXE2MEM_7_port, 
      NPC_EXE2MEM_6_port, NPC_EXE2MEM_5_port, NPC_EXE2MEM_4_port, 
      NPC_EXE2MEM_3_port, NPC_EXE2MEM_2_port, NPC_EXE2MEM_1_port, 
      NPC_EXE2MEM_0_port, ZOP_EXE2MEM, ALU_EXE2MEM_31_port, ALU_EXE2MEM_30_port
      , ALU_EXE2MEM_29_port, ALU_EXE2MEM_28_port, ALU_EXE2MEM_27_port, 
      ALU_EXE2MEM_26_port, ALU_EXE2MEM_25_port, ALU_EXE2MEM_24_port, 
      ALU_EXE2MEM_23_port, ALU_EXE2MEM_22_port, ALU_EXE2MEM_21_port, 
      ALU_EXE2MEM_20_port, ALU_EXE2MEM_19_port, ALU_EXE2MEM_18_port, 
      ALU_EXE2MEM_17_port, ALU_EXE2MEM_16_port, ALU_EXE2MEM_15_port, 
      ALU_EXE2MEM_14_port, ALU_EXE2MEM_13_port, ALU_EXE2MEM_12_port, 
      ALU_EXE2MEM_11_port, ALU_EXE2MEM_10_port, ALU_EXE2MEM_9_port, 
      ALU_EXE2MEM_8_port, ALU_EXE2MEM_7_port, ALU_EXE2MEM_6_port, 
      ALU_EXE2MEM_5_port, ALU_EXE2MEM_4_port, ALU_EXE2MEM_3_port, 
      ALU_EXE2MEM_2_port, ALU_EXE2MEM_1_port, ALU_EXE2MEM_0_port, 
      PAD_EXE2MEM_31_port, PAD_EXE2MEM_30_port, PAD_EXE2MEM_29_port, 
      PAD_EXE2MEM_28_port, PAD_EXE2MEM_27_port, PAD_EXE2MEM_26_port, 
      PAD_EXE2MEM_25_port, PAD_EXE2MEM_24_port, PAD_EXE2MEM_23_port, 
      PAD_EXE2MEM_22_port, PAD_EXE2MEM_21_port, PAD_EXE2MEM_20_port, 
      PAD_EXE2MEM_19_port, PAD_EXE2MEM_18_port, PAD_EXE2MEM_17_port, 
      PAD_EXE2MEM_16_port, PAD_EXE2MEM_15_port, PAD_EXE2MEM_14_port, 
      PAD_EXE2MEM_13_port, PAD_EXE2MEM_12_port, PAD_EXE2MEM_11_port, 
      PAD_EXE2MEM_10_port, PAD_EXE2MEM_9_port, PAD_EXE2MEM_8_port, 
      PAD_EXE2MEM_7_port, PAD_EXE2MEM_6_port, PAD_EXE2MEM_5_port, 
      PAD_EXE2MEM_4_port, PAD_EXE2MEM_3_port, PAD_EXE2MEM_2_port, 
      PAD_EXE2MEM_1_port, PAD_EXE2MEM_0_port, IR_EXE2MEM_4_port, 
      IR_EXE2MEM_3_port, IR_EXE2MEM_2_port, IR_EXE2MEM_1_port, 
      IR_EXE2MEM_0_port, IR_MEM2WB_4_port, IR_MEM2WB_3_port, IR_MEM2WB_2_port, 
      IR_MEM2WB_1_port, IR_MEM2WB_0_port, NPC_MEM2WB_31_port, 
      NPC_MEM2WB_30_port, NPC_MEM2WB_29_port, NPC_MEM2WB_28_port, 
      NPC_MEM2WB_27_port, NPC_MEM2WB_26_port, NPC_MEM2WB_25_port, 
      NPC_MEM2WB_24_port, NPC_MEM2WB_23_port, NPC_MEM2WB_22_port, 
      NPC_MEM2WB_21_port, NPC_MEM2WB_20_port, NPC_MEM2WB_19_port, 
      NPC_MEM2WB_18_port, NPC_MEM2WB_17_port, NPC_MEM2WB_16_port, 
      NPC_MEM2WB_15_port, NPC_MEM2WB_14_port, NPC_MEM2WB_13_port, 
      NPC_MEM2WB_12_port, NPC_MEM2WB_11_port, NPC_MEM2WB_10_port, 
      NPC_MEM2WB_9_port, NPC_MEM2WB_8_port, NPC_MEM2WB_7_port, 
      NPC_MEM2WB_6_port, NPC_MEM2WB_5_port, NPC_MEM2WB_4_port, 
      NPC_MEM2WB_3_port, NPC_MEM2WB_2_port, NPC_MEM2WB_1_port, 
      NPC_MEM2WB_0_port, ALU_MEM2WB_31_port, ALU_MEM2WB_30_port, 
      ALU_MEM2WB_29_port, ALU_MEM2WB_28_port, ALU_MEM2WB_27_port, 
      ALU_MEM2WB_26_port, ALU_MEM2WB_25_port, ALU_MEM2WB_24_port, 
      ALU_MEM2WB_23_port, ALU_MEM2WB_22_port, ALU_MEM2WB_21_port, 
      ALU_MEM2WB_20_port, ALU_MEM2WB_19_port, ALU_MEM2WB_18_port, 
      ALU_MEM2WB_17_port, ALU_MEM2WB_16_port, ALU_MEM2WB_15_port, 
      ALU_MEM2WB_14_port, ALU_MEM2WB_13_port, ALU_MEM2WB_12_port, 
      ALU_MEM2WB_11_port, ALU_MEM2WB_10_port, ALU_MEM2WB_9_port, 
      ALU_MEM2WB_8_port, ALU_MEM2WB_7_port, ALU_MEM2WB_6_port, 
      ALU_MEM2WB_5_port, ALU_MEM2WB_4_port, ALU_MEM2WB_3_port, 
      ALU_MEM2WB_2_port, ALU_MEM2WB_1_port, ALU_MEM2WB_0_port, 
      MEM_MEM2WB_31_port, MEM_MEM2WB_30_port, MEM_MEM2WB_29_port, 
      MEM_MEM2WB_28_port, MEM_MEM2WB_27_port, MEM_MEM2WB_26_port, 
      MEM_MEM2WB_25_port, MEM_MEM2WB_24_port, MEM_MEM2WB_23_port, 
      MEM_MEM2WB_22_port, MEM_MEM2WB_21_port, MEM_MEM2WB_20_port, 
      MEM_MEM2WB_19_port, MEM_MEM2WB_18_port, MEM_MEM2WB_17_port, 
      MEM_MEM2WB_16_port, MEM_MEM2WB_15_port, MEM_MEM2WB_14_port, 
      MEM_MEM2WB_13_port, MEM_MEM2WB_12_port, MEM_MEM2WB_11_port, 
      MEM_MEM2WB_10_port, MEM_MEM2WB_9_port, MEM_MEM2WB_8_port, 
      MEM_MEM2WB_7_port, MEM_MEM2WB_6_port, MEM_MEM2WB_5_port, 
      MEM_MEM2WB_4_port, MEM_MEM2WB_3_port, MEM_MEM2WB_2_port, 
      MEM_MEM2WB_1_port, MEM_MEM2WB_0_port, n_2208, n_2209, n_2210, n_2211 : 
      std_logic;

begin
   
   FETCH : IF_STAGE_N_BITS_DATA32_N_BYTES_INST4 port map( CLK => CLK, RST => 
                           RST, IF_LATCH_EN => IF_LATCH_EN, PC_LATCH_EN => 
                           PC_LATCH_EN, PC_IN(31) => PC_MEM2IF_31_port, 
                           PC_IN(30) => PC_MEM2IF_30_port, PC_IN(29) => 
                           PC_MEM2IF_29_port, PC_IN(28) => PC_MEM2IF_28_port, 
                           PC_IN(27) => PC_MEM2IF_27_port, PC_IN(26) => 
                           PC_MEM2IF_26_port, PC_IN(25) => PC_MEM2IF_25_port, 
                           PC_IN(24) => PC_MEM2IF_24_port, PC_IN(23) => 
                           PC_MEM2IF_23_port, PC_IN(22) => PC_MEM2IF_22_port, 
                           PC_IN(21) => PC_MEM2IF_21_port, PC_IN(20) => 
                           PC_MEM2IF_20_port, PC_IN(19) => PC_MEM2IF_19_port, 
                           PC_IN(18) => PC_MEM2IF_18_port, PC_IN(17) => 
                           PC_MEM2IF_17_port, PC_IN(16) => PC_MEM2IF_16_port, 
                           PC_IN(15) => PC_MEM2IF_15_port, PC_IN(14) => 
                           PC_MEM2IF_14_port, PC_IN(13) => PC_MEM2IF_13_port, 
                           PC_IN(12) => PC_MEM2IF_12_port, PC_IN(11) => 
                           PC_MEM2IF_11_port, PC_IN(10) => PC_MEM2IF_10_port, 
                           PC_IN(9) => PC_MEM2IF_9_port, PC_IN(8) => 
                           PC_MEM2IF_8_port, PC_IN(7) => PC_MEM2IF_7_port, 
                           PC_IN(6) => PC_MEM2IF_6_port, PC_IN(5) => 
                           PC_MEM2IF_5_port, PC_IN(4) => PC_MEM2IF_4_port, 
                           PC_IN(3) => PC_MEM2IF_3_port, PC_IN(2) => 
                           PC_MEM2IF_2_port, PC_IN(1) => PC_MEM2IF_1_port, 
                           PC_IN(0) => PC_MEM2IF_0_port, IR_IN(31) => IR_IN(31)
                           , IR_IN(30) => IR_IN(30), IR_IN(29) => IR_IN(29), 
                           IR_IN(28) => IR_IN(28), IR_IN(27) => IR_IN(27), 
                           IR_IN(26) => IR_IN(26), IR_IN(25) => IR_IN(25), 
                           IR_IN(24) => IR_IN(24), IR_IN(23) => IR_IN(23), 
                           IR_IN(22) => IR_IN(22), IR_IN(21) => IR_IN(21), 
                           IR_IN(20) => IR_IN(20), IR_IN(19) => IR_IN(19), 
                           IR_IN(18) => IR_IN(18), IR_IN(17) => IR_IN(17), 
                           IR_IN(16) => IR_IN(16), IR_IN(15) => IR_IN(15), 
                           IR_IN(14) => IR_IN(14), IR_IN(13) => IR_IN(13), 
                           IR_IN(12) => IR_IN(12), IR_IN(11) => IR_IN(11), 
                           IR_IN(10) => IR_IN(10), IR_IN(9) => IR_IN(9), 
                           IR_IN(8) => IR_IN(8), IR_IN(7) => IR_IN(7), IR_IN(6)
                           => IR_IN(6), IR_IN(5) => IR_IN(5), IR_IN(4) => 
                           IR_IN(4), IR_IN(3) => IR_IN(3), IR_IN(2) => IR_IN(2)
                           , IR_IN(1) => IR_IN(1), IR_IN(0) => IR_IN(0), 
                           PC_OUT(31) => PC_OUT(31), PC_OUT(30) => PC_OUT(30), 
                           PC_OUT(29) => PC_OUT(29), PC_OUT(28) => PC_OUT(28), 
                           PC_OUT(27) => PC_OUT(27), PC_OUT(26) => PC_OUT(26), 
                           PC_OUT(25) => PC_OUT(25), PC_OUT(24) => PC_OUT(24), 
                           PC_OUT(23) => PC_OUT(23), PC_OUT(22) => PC_OUT(22), 
                           PC_OUT(21) => PC_OUT(21), PC_OUT(20) => PC_OUT(20), 
                           PC_OUT(19) => PC_OUT(19), PC_OUT(18) => PC_OUT(18), 
                           PC_OUT(17) => PC_OUT(17), PC_OUT(16) => PC_OUT(16), 
                           PC_OUT(15) => PC_OUT(15), PC_OUT(14) => PC_OUT(14), 
                           PC_OUT(13) => PC_OUT(13), PC_OUT(12) => PC_OUT(12), 
                           PC_OUT(11) => PC_OUT(11), PC_OUT(10) => PC_OUT(10), 
                           PC_OUT(9) => PC_OUT(9), PC_OUT(8) => PC_OUT(8), 
                           PC_OUT(7) => PC_OUT(7), PC_OUT(6) => PC_OUT(6), 
                           PC_OUT(5) => PC_OUT(5), PC_OUT(4) => PC_OUT(4), 
                           PC_OUT(3) => PC_OUT(3), PC_OUT(2) => PC_OUT(2), 
                           PC_OUT(1) => PC_OUT(1), PC_OUT(0) => PC_OUT(0), 
                           IR_OUT(31) => IR_IF2ID_31_port, IR_OUT(30) => 
                           IR_IF2ID_30_port, IR_OUT(29) => IR_IF2ID_29_port, 
                           IR_OUT(28) => IR_IF2ID_28_port, IR_OUT(27) => 
                           IR_IF2ID_27_port, IR_OUT(26) => IR_IF2ID_26_port, 
                           IR_OUT(25) => IR_IF2ID_25_port, IR_OUT(24) => 
                           IR_IF2ID_24_port, IR_OUT(23) => IR_IF2ID_23_port, 
                           IR_OUT(22) => IR_IF2ID_22_port, IR_OUT(21) => 
                           IR_IF2ID_21_port, IR_OUT(20) => IR_IF2ID_20_port, 
                           IR_OUT(19) => IR_IF2ID_19_port, IR_OUT(18) => 
                           IR_IF2ID_18_port, IR_OUT(17) => IR_IF2ID_17_port, 
                           IR_OUT(16) => IR_IF2ID_16_port, IR_OUT(15) => 
                           IR_IF2ID_15_port, IR_OUT(14) => IR_IF2ID_14_port, 
                           IR_OUT(13) => IR_IF2ID_13_port, IR_OUT(12) => 
                           IR_IF2ID_12_port, IR_OUT(11) => IR_IF2ID_11_port, 
                           IR_OUT(10) => IR_IF2ID_10_port, IR_OUT(9) => 
                           IR_IF2ID_9_port, IR_OUT(8) => IR_IF2ID_8_port, 
                           IR_OUT(7) => IR_IF2ID_7_port, IR_OUT(6) => 
                           IR_IF2ID_6_port, IR_OUT(5) => IR_IF2ID_5_port, 
                           IR_OUT(4) => IR_IF2ID_4_port, IR_OUT(3) => 
                           IR_IF2ID_3_port, IR_OUT(2) => IR_IF2ID_2_port, 
                           IR_OUT(1) => IR_IF2ID_1_port, IR_OUT(0) => 
                           IR_IF2ID_0_port, NPC_OUT(31) => 
                           NPC_IF2ID_MEM_31_port, NPC_OUT(30) => 
                           NPC_IF2ID_MEM_30_port, NPC_OUT(29) => 
                           NPC_IF2ID_MEM_29_port, NPC_OUT(28) => 
                           NPC_IF2ID_MEM_28_port, NPC_OUT(27) => 
                           NPC_IF2ID_MEM_27_port, NPC_OUT(26) => 
                           NPC_IF2ID_MEM_26_port, NPC_OUT(25) => 
                           NPC_IF2ID_MEM_25_port, NPC_OUT(24) => 
                           NPC_IF2ID_MEM_24_port, NPC_OUT(23) => 
                           NPC_IF2ID_MEM_23_port, NPC_OUT(22) => 
                           NPC_IF2ID_MEM_22_port, NPC_OUT(21) => 
                           NPC_IF2ID_MEM_21_port, NPC_OUT(20) => 
                           NPC_IF2ID_MEM_20_port, NPC_OUT(19) => 
                           NPC_IF2ID_MEM_19_port, NPC_OUT(18) => 
                           NPC_IF2ID_MEM_18_port, NPC_OUT(17) => 
                           NPC_IF2ID_MEM_17_port, NPC_OUT(16) => 
                           NPC_IF2ID_MEM_16_port, NPC_OUT(15) => 
                           NPC_IF2ID_MEM_15_port, NPC_OUT(14) => 
                           NPC_IF2ID_MEM_14_port, NPC_OUT(13) => 
                           NPC_IF2ID_MEM_13_port, NPC_OUT(12) => 
                           NPC_IF2ID_MEM_12_port, NPC_OUT(11) => 
                           NPC_IF2ID_MEM_11_port, NPC_OUT(10) => 
                           NPC_IF2ID_MEM_10_port, NPC_OUT(9) => 
                           NPC_IF2ID_MEM_9_port, NPC_OUT(8) => 
                           NPC_IF2ID_MEM_8_port, NPC_OUT(7) => 
                           NPC_IF2ID_MEM_7_port, NPC_OUT(6) => 
                           NPC_IF2ID_MEM_6_port, NPC_OUT(5) => 
                           NPC_IF2ID_MEM_5_port, NPC_OUT(4) => 
                           NPC_IF2ID_MEM_4_port, NPC_OUT(3) => 
                           NPC_IF2ID_MEM_3_port, NPC_OUT(2) => 
                           NPC_IF2ID_MEM_2_port, NPC_OUT(1) => 
                           NPC_IF2ID_MEM_1_port, NPC_OUT(0) => 
                           NPC_IF2ID_MEM_0_port);
   DECODE : 
                           ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 
                           port map( CLK => CLK, RST => RST, JAL_MUX_SEL => 
                           JAL_MUX_SEL, DEC_OUTREG_EN => DEC_OUTREG_EN, 
                           IS_I_TYPE => IS_I_TYPE, RD1_EN => RD1_EN, RD2_EN => 
                           RD2_EN, WR_EN => WR_EN, ZERO_PADDING2 => 
                           ZERO_PADDING2, I_CODE(31) => IR_IF2ID_31_port, 
                           I_CODE(30) => IR_IF2ID_30_port, I_CODE(29) => 
                           IR_IF2ID_29_port, I_CODE(28) => IR_IF2ID_28_port, 
                           I_CODE(27) => IR_IF2ID_27_port, I_CODE(26) => 
                           IR_IF2ID_26_port, I_CODE(25) => IR_IF2ID_25_port, 
                           I_CODE(24) => IR_IF2ID_24_port, I_CODE(23) => 
                           IR_IF2ID_23_port, I_CODE(22) => IR_IF2ID_22_port, 
                           I_CODE(21) => IR_IF2ID_21_port, I_CODE(20) => 
                           IR_IF2ID_20_port, I_CODE(19) => IR_IF2ID_19_port, 
                           I_CODE(18) => IR_IF2ID_18_port, I_CODE(17) => 
                           IR_IF2ID_17_port, I_CODE(16) => IR_IF2ID_16_port, 
                           I_CODE(15) => IR_IF2ID_15_port, I_CODE(14) => 
                           IR_IF2ID_14_port, I_CODE(13) => IR_IF2ID_13_port, 
                           I_CODE(12) => IR_IF2ID_12_port, I_CODE(11) => 
                           IR_IF2ID_11_port, I_CODE(10) => IR_IF2ID_10_port, 
                           I_CODE(9) => IR_IF2ID_9_port, I_CODE(8) => 
                           IR_IF2ID_8_port, I_CODE(7) => IR_IF2ID_7_port, 
                           I_CODE(6) => IR_IF2ID_6_port, I_CODE(5) => 
                           IR_IF2ID_5_port, I_CODE(4) => IR_IF2ID_4_port, 
                           I_CODE(3) => IR_IF2ID_3_port, I_CODE(2) => 
                           IR_IF2ID_2_port, I_CODE(1) => IR_IF2ID_1_port, 
                           I_CODE(0) => IR_IF2ID_0_port, NPC1_IN(31) => 
                           NPC_IF2ID_MEM_31_port, NPC1_IN(30) => 
                           NPC_IF2ID_MEM_30_port, NPC1_IN(29) => 
                           NPC_IF2ID_MEM_29_port, NPC1_IN(28) => 
                           NPC_IF2ID_MEM_28_port, NPC1_IN(27) => 
                           NPC_IF2ID_MEM_27_port, NPC1_IN(26) => 
                           NPC_IF2ID_MEM_26_port, NPC1_IN(25) => 
                           NPC_IF2ID_MEM_25_port, NPC1_IN(24) => 
                           NPC_IF2ID_MEM_24_port, NPC1_IN(23) => 
                           NPC_IF2ID_MEM_23_port, NPC1_IN(22) => 
                           NPC_IF2ID_MEM_22_port, NPC1_IN(21) => 
                           NPC_IF2ID_MEM_21_port, NPC1_IN(20) => 
                           NPC_IF2ID_MEM_20_port, NPC1_IN(19) => 
                           NPC_IF2ID_MEM_19_port, NPC1_IN(18) => 
                           NPC_IF2ID_MEM_18_port, NPC1_IN(17) => 
                           NPC_IF2ID_MEM_17_port, NPC1_IN(16) => 
                           NPC_IF2ID_MEM_16_port, NPC1_IN(15) => 
                           NPC_IF2ID_MEM_15_port, NPC1_IN(14) => 
                           NPC_IF2ID_MEM_14_port, NPC1_IN(13) => 
                           NPC_IF2ID_MEM_13_port, NPC1_IN(12) => 
                           NPC_IF2ID_MEM_12_port, NPC1_IN(11) => 
                           NPC_IF2ID_MEM_11_port, NPC1_IN(10) => 
                           NPC_IF2ID_MEM_10_port, NPC1_IN(9) => 
                           NPC_IF2ID_MEM_9_port, NPC1_IN(8) => 
                           NPC_IF2ID_MEM_8_port, NPC1_IN(7) => 
                           NPC_IF2ID_MEM_7_port, NPC1_IN(6) => 
                           NPC_IF2ID_MEM_6_port, NPC1_IN(5) => 
                           NPC_IF2ID_MEM_5_port, NPC1_IN(4) => 
                           NPC_IF2ID_MEM_4_port, NPC1_IN(3) => 
                           NPC_IF2ID_MEM_3_port, NPC1_IN(2) => 
                           NPC_IF2ID_MEM_2_port, NPC1_IN(1) => 
                           NPC_IF2ID_MEM_1_port, NPC1_IN(0) => 
                           NPC_IF2ID_MEM_0_port, DATA_IN(31) => 
                           WRT_WB2ID_31_port, DATA_IN(30) => WRT_WB2ID_30_port,
                           DATA_IN(29) => WRT_WB2ID_29_port, DATA_IN(28) => 
                           WRT_WB2ID_28_port, DATA_IN(27) => WRT_WB2ID_27_port,
                           DATA_IN(26) => WRT_WB2ID_26_port, DATA_IN(25) => 
                           WRT_WB2ID_25_port, DATA_IN(24) => WRT_WB2ID_24_port,
                           DATA_IN(23) => WRT_WB2ID_23_port, DATA_IN(22) => 
                           WRT_WB2ID_22_port, DATA_IN(21) => WRT_WB2ID_21_port,
                           DATA_IN(20) => WRT_WB2ID_20_port, DATA_IN(19) => 
                           WRT_WB2ID_19_port, DATA_IN(18) => WRT_WB2ID_18_port,
                           DATA_IN(17) => WRT_WB2ID_17_port, DATA_IN(16) => 
                           WRT_WB2ID_16_port, DATA_IN(15) => WRT_WB2ID_15_port,
                           DATA_IN(14) => WRT_WB2ID_14_port, DATA_IN(13) => 
                           WRT_WB2ID_13_port, DATA_IN(12) => WRT_WB2ID_12_port,
                           DATA_IN(11) => WRT_WB2ID_11_port, DATA_IN(10) => 
                           WRT_WB2ID_10_port, DATA_IN(9) => WRT_WB2ID_9_port, 
                           DATA_IN(8) => WRT_WB2ID_8_port, DATA_IN(7) => 
                           WRT_WB2ID_7_port, DATA_IN(6) => WRT_WB2ID_6_port, 
                           DATA_IN(5) => WRT_WB2ID_5_port, DATA_IN(4) => 
                           WRT_WB2ID_4_port, DATA_IN(3) => WRT_WB2ID_3_port, 
                           DATA_IN(2) => WRT_WB2ID_2_port, DATA_IN(1) => 
                           WRT_WB2ID_1_port, DATA_IN(0) => WRT_WB2ID_0_port, 
                           WR_ADDR_IN(4) => IR_WB2ID_4_port, WR_ADDR_IN(3) => 
                           IR_WB2ID_3_port, WR_ADDR_IN(2) => IR_WB2ID_2_port, 
                           WR_ADDR_IN(1) => IR_WB2ID_1_port, WR_ADDR_IN(0) => 
                           IR_WB2ID_0_port, REGA_OUT(31) => A_ID2EXE_31_port, 
                           REGA_OUT(30) => A_ID2EXE_30_port, REGA_OUT(29) => 
                           A_ID2EXE_29_port, REGA_OUT(28) => A_ID2EXE_28_port, 
                           REGA_OUT(27) => A_ID2EXE_27_port, REGA_OUT(26) => 
                           A_ID2EXE_26_port, REGA_OUT(25) => A_ID2EXE_25_port, 
                           REGA_OUT(24) => A_ID2EXE_24_port, REGA_OUT(23) => 
                           A_ID2EXE_23_port, REGA_OUT(22) => A_ID2EXE_22_port, 
                           REGA_OUT(21) => A_ID2EXE_21_port, REGA_OUT(20) => 
                           A_ID2EXE_20_port, REGA_OUT(19) => A_ID2EXE_19_port, 
                           REGA_OUT(18) => A_ID2EXE_18_port, REGA_OUT(17) => 
                           A_ID2EXE_17_port, REGA_OUT(16) => A_ID2EXE_16_port, 
                           REGA_OUT(15) => A_ID2EXE_15_port, REGA_OUT(14) => 
                           A_ID2EXE_14_port, REGA_OUT(13) => A_ID2EXE_13_port, 
                           REGA_OUT(12) => A_ID2EXE_12_port, REGA_OUT(11) => 
                           A_ID2EXE_11_port, REGA_OUT(10) => A_ID2EXE_10_port, 
                           REGA_OUT(9) => A_ID2EXE_9_port, REGA_OUT(8) => 
                           A_ID2EXE_8_port, REGA_OUT(7) => A_ID2EXE_7_port, 
                           REGA_OUT(6) => A_ID2EXE_6_port, REGA_OUT(5) => 
                           A_ID2EXE_5_port, REGA_OUT(4) => A_ID2EXE_4_port, 
                           REGA_OUT(3) => A_ID2EXE_3_port, REGA_OUT(2) => 
                           A_ID2EXE_2_port, REGA_OUT(1) => A_ID2EXE_1_port, 
                           REGA_OUT(0) => A_ID2EXE_0_port, REGB_OUT(31) => 
                           B_ID2EXE_31_port, REGB_OUT(30) => B_ID2EXE_30_port, 
                           REGB_OUT(29) => B_ID2EXE_29_port, REGB_OUT(28) => 
                           B_ID2EXE_28_port, REGB_OUT(27) => B_ID2EXE_27_port, 
                           REGB_OUT(26) => B_ID2EXE_26_port, REGB_OUT(25) => 
                           B_ID2EXE_25_port, REGB_OUT(24) => B_ID2EXE_24_port, 
                           REGB_OUT(23) => B_ID2EXE_23_port, REGB_OUT(22) => 
                           B_ID2EXE_22_port, REGB_OUT(21) => B_ID2EXE_21_port, 
                           REGB_OUT(20) => B_ID2EXE_20_port, REGB_OUT(19) => 
                           B_ID2EXE_19_port, REGB_OUT(18) => B_ID2EXE_18_port, 
                           REGB_OUT(17) => B_ID2EXE_17_port, REGB_OUT(16) => 
                           B_ID2EXE_16_port, REGB_OUT(15) => B_ID2EXE_15_port, 
                           REGB_OUT(14) => B_ID2EXE_14_port, REGB_OUT(13) => 
                           B_ID2EXE_13_port, REGB_OUT(12) => B_ID2EXE_12_port, 
                           REGB_OUT(11) => B_ID2EXE_11_port, REGB_OUT(10) => 
                           B_ID2EXE_10_port, REGB_OUT(9) => B_ID2EXE_9_port, 
                           REGB_OUT(8) => B_ID2EXE_8_port, REGB_OUT(7) => 
                           B_ID2EXE_7_port, REGB_OUT(6) => B_ID2EXE_6_port, 
                           REGB_OUT(5) => B_ID2EXE_5_port, REGB_OUT(4) => 
                           B_ID2EXE_4_port, REGB_OUT(3) => B_ID2EXE_3_port, 
                           REGB_OUT(2) => B_ID2EXE_2_port, REGB_OUT(1) => 
                           B_ID2EXE_1_port, REGB_OUT(0) => B_ID2EXE_0_port, 
                           REGIMM_OUT(31) => IMM_ID2EXE_31_port, REGIMM_OUT(30)
                           => IMM_ID2EXE_30_port, REGIMM_OUT(29) => 
                           IMM_ID2EXE_29_port, REGIMM_OUT(28) => 
                           IMM_ID2EXE_28_port, REGIMM_OUT(27) => 
                           IMM_ID2EXE_27_port, REGIMM_OUT(26) => 
                           IMM_ID2EXE_26_port, REGIMM_OUT(25) => 
                           IMM_ID2EXE_25_port, REGIMM_OUT(24) => 
                           IMM_ID2EXE_24_port, REGIMM_OUT(23) => 
                           IMM_ID2EXE_23_port, REGIMM_OUT(22) => 
                           IMM_ID2EXE_22_port, REGIMM_OUT(21) => 
                           IMM_ID2EXE_21_port, REGIMM_OUT(20) => 
                           IMM_ID2EXE_20_port, REGIMM_OUT(19) => 
                           IMM_ID2EXE_19_port, REGIMM_OUT(18) => 
                           IMM_ID2EXE_18_port, REGIMM_OUT(17) => 
                           IMM_ID2EXE_17_port, REGIMM_OUT(16) => 
                           IMM_ID2EXE_16_port, REGIMM_OUT(15) => 
                           IMM_ID2EXE_15_port, REGIMM_OUT(14) => 
                           IMM_ID2EXE_14_port, REGIMM_OUT(13) => 
                           IMM_ID2EXE_13_port, REGIMM_OUT(12) => 
                           IMM_ID2EXE_12_port, REGIMM_OUT(11) => 
                           IMM_ID2EXE_11_port, REGIMM_OUT(10) => 
                           IMM_ID2EXE_10_port, REGIMM_OUT(9) => 
                           IMM_ID2EXE_9_port, REGIMM_OUT(8) => 
                           IMM_ID2EXE_8_port, REGIMM_OUT(7) => 
                           IMM_ID2EXE_7_port, REGIMM_OUT(6) => 
                           IMM_ID2EXE_6_port, REGIMM_OUT(5) => 
                           IMM_ID2EXE_5_port, REGIMM_OUT(4) => 
                           IMM_ID2EXE_4_port, REGIMM_OUT(3) => 
                           IMM_ID2EXE_3_port, REGIMM_OUT(2) => 
                           IMM_ID2EXE_2_port, REGIMM_OUT(1) => 
                           IMM_ID2EXE_1_port, REGIMM_OUT(0) => 
                           IMM_ID2EXE_0_port, WR_ADDR_OUT(4) => 
                           IR_ID2EXE_4_port, WR_ADDR_OUT(3) => IR_ID2EXE_3_port
                           , WR_ADDR_OUT(2) => IR_ID2EXE_2_port, WR_ADDR_OUT(1)
                           => IR_ID2EXE_1_port, WR_ADDR_OUT(0) => 
                           IR_ID2EXE_0_port, NPC1_OUT(31) => NPC_ID2EXE_31_port
                           , NPC1_OUT(30) => NPC_ID2EXE_30_port, NPC1_OUT(29) 
                           => NPC_ID2EXE_29_port, NPC1_OUT(28) => 
                           NPC_ID2EXE_28_port, NPC1_OUT(27) => 
                           NPC_ID2EXE_27_port, NPC1_OUT(26) => 
                           NPC_ID2EXE_26_port, NPC1_OUT(25) => 
                           NPC_ID2EXE_25_port, NPC1_OUT(24) => 
                           NPC_ID2EXE_24_port, NPC1_OUT(23) => 
                           NPC_ID2EXE_23_port, NPC1_OUT(22) => 
                           NPC_ID2EXE_22_port, NPC1_OUT(21) => 
                           NPC_ID2EXE_21_port, NPC1_OUT(20) => 
                           NPC_ID2EXE_20_port, NPC1_OUT(19) => 
                           NPC_ID2EXE_19_port, NPC1_OUT(18) => 
                           NPC_ID2EXE_18_port, NPC1_OUT(17) => 
                           NPC_ID2EXE_17_port, NPC1_OUT(16) => 
                           NPC_ID2EXE_16_port, NPC1_OUT(15) => 
                           NPC_ID2EXE_15_port, NPC1_OUT(14) => 
                           NPC_ID2EXE_14_port, NPC1_OUT(13) => 
                           NPC_ID2EXE_13_port, NPC1_OUT(12) => 
                           NPC_ID2EXE_12_port, NPC1_OUT(11) => 
                           NPC_ID2EXE_11_port, NPC1_OUT(10) => 
                           NPC_ID2EXE_10_port, NPC1_OUT(9) => NPC_ID2EXE_9_port
                           , NPC1_OUT(8) => NPC_ID2EXE_8_port, NPC1_OUT(7) => 
                           NPC_ID2EXE_7_port, NPC1_OUT(6) => NPC_ID2EXE_6_port,
                           NPC1_OUT(5) => NPC_ID2EXE_5_port, NPC1_OUT(4) => 
                           NPC_ID2EXE_4_port, NPC1_OUT(3) => NPC_ID2EXE_3_port,
                           NPC1_OUT(2) => NPC_ID2EXE_2_port, NPC1_OUT(1) => 
                           NPC_ID2EXE_1_port, NPC1_OUT(0) => NPC_ID2EXE_0_port)
                           ;
   EXECUTE : EXE_STAGE_N_BITS_DATA32_RF_ADDR5 port map( CLK => CLK, RST => RST,
                           MUXA_SEL => MUXA_SEL, MUXB_SEL => MUXB_SEL, 
                           EXE_OUTREG_EN => EXE_OUTREG_EN, EQ_COND => EQ_COND, 
                           JUMP_EN => JUMP_EN, ALU_OPCODE(0) => ALU_OPCODE(0), 
                           ALU_OPCODE(1) => ALU_OPCODE(1), ALU_OPCODE(2) => 
                           ALU_OPCODE(2), ALU_OPCODE(3) => ALU_OPCODE(3), 
                           ALU_OPCODE(4) => ALU_OPCODE(4), ALU_OPCODE(5) => 
                           ALU_OPCODE(5), ALU_OPCODE(6) => ALU_OPCODE(6), 
                           NPC2_IN(31) => NPC_ID2EXE_31_port, NPC2_IN(30) => 
                           NPC_ID2EXE_30_port, NPC2_IN(29) => 
                           NPC_ID2EXE_29_port, NPC2_IN(28) => 
                           NPC_ID2EXE_28_port, NPC2_IN(27) => 
                           NPC_ID2EXE_27_port, NPC2_IN(26) => 
                           NPC_ID2EXE_26_port, NPC2_IN(25) => 
                           NPC_ID2EXE_25_port, NPC2_IN(24) => 
                           NPC_ID2EXE_24_port, NPC2_IN(23) => 
                           NPC_ID2EXE_23_port, NPC2_IN(22) => 
                           NPC_ID2EXE_22_port, NPC2_IN(21) => 
                           NPC_ID2EXE_21_port, NPC2_IN(20) => 
                           NPC_ID2EXE_20_port, NPC2_IN(19) => 
                           NPC_ID2EXE_19_port, NPC2_IN(18) => 
                           NPC_ID2EXE_18_port, NPC2_IN(17) => 
                           NPC_ID2EXE_17_port, NPC2_IN(16) => 
                           NPC_ID2EXE_16_port, NPC2_IN(15) => 
                           NPC_ID2EXE_15_port, NPC2_IN(14) => 
                           NPC_ID2EXE_14_port, NPC2_IN(13) => 
                           NPC_ID2EXE_13_port, NPC2_IN(12) => 
                           NPC_ID2EXE_12_port, NPC2_IN(11) => 
                           NPC_ID2EXE_11_port, NPC2_IN(10) => 
                           NPC_ID2EXE_10_port, NPC2_IN(9) => NPC_ID2EXE_9_port,
                           NPC2_IN(8) => NPC_ID2EXE_8_port, NPC2_IN(7) => 
                           NPC_ID2EXE_7_port, NPC2_IN(6) => NPC_ID2EXE_6_port, 
                           NPC2_IN(5) => NPC_ID2EXE_5_port, NPC2_IN(4) => 
                           NPC_ID2EXE_4_port, NPC2_IN(3) => NPC_ID2EXE_3_port, 
                           NPC2_IN(2) => NPC_ID2EXE_2_port, NPC2_IN(1) => 
                           NPC_ID2EXE_1_port, NPC2_IN(0) => NPC_ID2EXE_0_port, 
                           NPC1_MUXA_IN(31) => NPC_ID2EXE_31_port, 
                           NPC1_MUXA_IN(30) => NPC_ID2EXE_30_port, 
                           NPC1_MUXA_IN(29) => NPC_ID2EXE_29_port, 
                           NPC1_MUXA_IN(28) => NPC_ID2EXE_28_port, 
                           NPC1_MUXA_IN(27) => NPC_ID2EXE_27_port, 
                           NPC1_MUXA_IN(26) => NPC_ID2EXE_26_port, 
                           NPC1_MUXA_IN(25) => NPC_ID2EXE_25_port, 
                           NPC1_MUXA_IN(24) => NPC_ID2EXE_24_port, 
                           NPC1_MUXA_IN(23) => NPC_ID2EXE_23_port, 
                           NPC1_MUXA_IN(22) => NPC_ID2EXE_22_port, 
                           NPC1_MUXA_IN(21) => NPC_ID2EXE_21_port, 
                           NPC1_MUXA_IN(20) => NPC_ID2EXE_20_port, 
                           NPC1_MUXA_IN(19) => NPC_ID2EXE_19_port, 
                           NPC1_MUXA_IN(18) => NPC_ID2EXE_18_port, 
                           NPC1_MUXA_IN(17) => NPC_ID2EXE_17_port, 
                           NPC1_MUXA_IN(16) => NPC_ID2EXE_16_port, 
                           NPC1_MUXA_IN(15) => NPC_ID2EXE_15_port, 
                           NPC1_MUXA_IN(14) => NPC_ID2EXE_14_port, 
                           NPC1_MUXA_IN(13) => NPC_ID2EXE_13_port, 
                           NPC1_MUXA_IN(12) => NPC_ID2EXE_12_port, 
                           NPC1_MUXA_IN(11) => NPC_ID2EXE_11_port, 
                           NPC1_MUXA_IN(10) => NPC_ID2EXE_10_port, 
                           NPC1_MUXA_IN(9) => NPC_ID2EXE_9_port, 
                           NPC1_MUXA_IN(8) => NPC_ID2EXE_8_port, 
                           NPC1_MUXA_IN(7) => NPC_ID2EXE_7_port, 
                           NPC1_MUXA_IN(6) => NPC_ID2EXE_6_port, 
                           NPC1_MUXA_IN(5) => NPC_ID2EXE_5_port, 
                           NPC1_MUXA_IN(4) => NPC_ID2EXE_4_port, 
                           NPC1_MUXA_IN(3) => NPC_ID2EXE_3_port, 
                           NPC1_MUXA_IN(2) => NPC_ID2EXE_2_port, 
                           NPC1_MUXA_IN(1) => NPC_ID2EXE_1_port, 
                           NPC1_MUXA_IN(0) => NPC_ID2EXE_0_port, 
                           REGA_MUXA_IN(31) => A_ID2EXE_31_port, 
                           REGA_MUXA_IN(30) => A_ID2EXE_30_port, 
                           REGA_MUXA_IN(29) => A_ID2EXE_29_port, 
                           REGA_MUXA_IN(28) => A_ID2EXE_28_port, 
                           REGA_MUXA_IN(27) => A_ID2EXE_27_port, 
                           REGA_MUXA_IN(26) => A_ID2EXE_26_port, 
                           REGA_MUXA_IN(25) => A_ID2EXE_25_port, 
                           REGA_MUXA_IN(24) => A_ID2EXE_24_port, 
                           REGA_MUXA_IN(23) => A_ID2EXE_23_port, 
                           REGA_MUXA_IN(22) => A_ID2EXE_22_port, 
                           REGA_MUXA_IN(21) => A_ID2EXE_21_port, 
                           REGA_MUXA_IN(20) => A_ID2EXE_20_port, 
                           REGA_MUXA_IN(19) => A_ID2EXE_19_port, 
                           REGA_MUXA_IN(18) => A_ID2EXE_18_port, 
                           REGA_MUXA_IN(17) => A_ID2EXE_17_port, 
                           REGA_MUXA_IN(16) => A_ID2EXE_16_port, 
                           REGA_MUXA_IN(15) => A_ID2EXE_15_port, 
                           REGA_MUXA_IN(14) => A_ID2EXE_14_port, 
                           REGA_MUXA_IN(13) => A_ID2EXE_13_port, 
                           REGA_MUXA_IN(12) => A_ID2EXE_12_port, 
                           REGA_MUXA_IN(11) => A_ID2EXE_11_port, 
                           REGA_MUXA_IN(10) => A_ID2EXE_10_port, 
                           REGA_MUXA_IN(9) => A_ID2EXE_9_port, REGA_MUXA_IN(8) 
                           => A_ID2EXE_8_port, REGA_MUXA_IN(7) => 
                           A_ID2EXE_7_port, REGA_MUXA_IN(6) => A_ID2EXE_6_port,
                           REGA_MUXA_IN(5) => A_ID2EXE_5_port, REGA_MUXA_IN(4) 
                           => A_ID2EXE_4_port, REGA_MUXA_IN(3) => 
                           A_ID2EXE_3_port, REGA_MUXA_IN(2) => A_ID2EXE_2_port,
                           REGA_MUXA_IN(1) => A_ID2EXE_1_port, REGA_MUXA_IN(0) 
                           => A_ID2EXE_0_port, REGB_MUXB_IN(31) => 
                           B_ID2EXE_31_port, REGB_MUXB_IN(30) => 
                           B_ID2EXE_30_port, REGB_MUXB_IN(29) => 
                           B_ID2EXE_29_port, REGB_MUXB_IN(28) => 
                           B_ID2EXE_28_port, REGB_MUXB_IN(27) => 
                           B_ID2EXE_27_port, REGB_MUXB_IN(26) => 
                           B_ID2EXE_26_port, REGB_MUXB_IN(25) => 
                           B_ID2EXE_25_port, REGB_MUXB_IN(24) => 
                           B_ID2EXE_24_port, REGB_MUXB_IN(23) => 
                           B_ID2EXE_23_port, REGB_MUXB_IN(22) => 
                           B_ID2EXE_22_port, REGB_MUXB_IN(21) => 
                           B_ID2EXE_21_port, REGB_MUXB_IN(20) => 
                           B_ID2EXE_20_port, REGB_MUXB_IN(19) => 
                           B_ID2EXE_19_port, REGB_MUXB_IN(18) => 
                           B_ID2EXE_18_port, REGB_MUXB_IN(17) => 
                           B_ID2EXE_17_port, REGB_MUXB_IN(16) => 
                           B_ID2EXE_16_port, REGB_MUXB_IN(15) => 
                           B_ID2EXE_15_port, REGB_MUXB_IN(14) => 
                           B_ID2EXE_14_port, REGB_MUXB_IN(13) => 
                           B_ID2EXE_13_port, REGB_MUXB_IN(12) => 
                           B_ID2EXE_12_port, REGB_MUXB_IN(11) => 
                           B_ID2EXE_11_port, REGB_MUXB_IN(10) => 
                           B_ID2EXE_10_port, REGB_MUXB_IN(9) => B_ID2EXE_9_port
                           , REGB_MUXB_IN(8) => B_ID2EXE_8_port, 
                           REGB_MUXB_IN(7) => B_ID2EXE_7_port, REGB_MUXB_IN(6) 
                           => B_ID2EXE_6_port, REGB_MUXB_IN(5) => 
                           B_ID2EXE_5_port, REGB_MUXB_IN(4) => B_ID2EXE_4_port,
                           REGB_MUXB_IN(3) => B_ID2EXE_3_port, REGB_MUXB_IN(2) 
                           => B_ID2EXE_2_port, REGB_MUXB_IN(1) => 
                           B_ID2EXE_1_port, REGB_MUXB_IN(0) => B_ID2EXE_0_port,
                           IMM_MUXB_IN(31) => IMM_ID2EXE_31_port, 
                           IMM_MUXB_IN(30) => IMM_ID2EXE_30_port, 
                           IMM_MUXB_IN(29) => IMM_ID2EXE_29_port, 
                           IMM_MUXB_IN(28) => IMM_ID2EXE_28_port, 
                           IMM_MUXB_IN(27) => IMM_ID2EXE_27_port, 
                           IMM_MUXB_IN(26) => IMM_ID2EXE_26_port, 
                           IMM_MUXB_IN(25) => IMM_ID2EXE_25_port, 
                           IMM_MUXB_IN(24) => IMM_ID2EXE_24_port, 
                           IMM_MUXB_IN(23) => IMM_ID2EXE_23_port, 
                           IMM_MUXB_IN(22) => IMM_ID2EXE_22_port, 
                           IMM_MUXB_IN(21) => IMM_ID2EXE_21_port, 
                           IMM_MUXB_IN(20) => IMM_ID2EXE_20_port, 
                           IMM_MUXB_IN(19) => IMM_ID2EXE_19_port, 
                           IMM_MUXB_IN(18) => IMM_ID2EXE_18_port, 
                           IMM_MUXB_IN(17) => IMM_ID2EXE_17_port, 
                           IMM_MUXB_IN(16) => IMM_ID2EXE_16_port, 
                           IMM_MUXB_IN(15) => IMM_ID2EXE_15_port, 
                           IMM_MUXB_IN(14) => IMM_ID2EXE_14_port, 
                           IMM_MUXB_IN(13) => IMM_ID2EXE_13_port, 
                           IMM_MUXB_IN(12) => IMM_ID2EXE_12_port, 
                           IMM_MUXB_IN(11) => IMM_ID2EXE_11_port, 
                           IMM_MUXB_IN(10) => IMM_ID2EXE_10_port, 
                           IMM_MUXB_IN(9) => IMM_ID2EXE_9_port, IMM_MUXB_IN(8) 
                           => IMM_ID2EXE_8_port, IMM_MUXB_IN(7) => 
                           IMM_ID2EXE_7_port, IMM_MUXB_IN(6) => 
                           IMM_ID2EXE_6_port, IMM_MUXB_IN(5) => 
                           IMM_ID2EXE_5_port, IMM_MUXB_IN(4) => 
                           IMM_ID2EXE_4_port, IMM_MUXB_IN(3) => 
                           IMM_ID2EXE_3_port, IMM_MUXB_IN(2) => 
                           IMM_ID2EXE_2_port, IMM_MUXB_IN(1) => 
                           IMM_ID2EXE_1_port, IMM_MUXB_IN(0) => 
                           IMM_ID2EXE_0_port, PAD_IN(31) => B_ID2EXE_31_port, 
                           PAD_IN(30) => B_ID2EXE_30_port, PAD_IN(29) => 
                           B_ID2EXE_29_port, PAD_IN(28) => B_ID2EXE_28_port, 
                           PAD_IN(27) => B_ID2EXE_27_port, PAD_IN(26) => 
                           B_ID2EXE_26_port, PAD_IN(25) => B_ID2EXE_25_port, 
                           PAD_IN(24) => B_ID2EXE_24_port, PAD_IN(23) => 
                           B_ID2EXE_23_port, PAD_IN(22) => B_ID2EXE_22_port, 
                           PAD_IN(21) => B_ID2EXE_21_port, PAD_IN(20) => 
                           B_ID2EXE_20_port, PAD_IN(19) => B_ID2EXE_19_port, 
                           PAD_IN(18) => B_ID2EXE_18_port, PAD_IN(17) => 
                           B_ID2EXE_17_port, PAD_IN(16) => B_ID2EXE_16_port, 
                           PAD_IN(15) => B_ID2EXE_15_port, PAD_IN(14) => 
                           B_ID2EXE_14_port, PAD_IN(13) => B_ID2EXE_13_port, 
                           PAD_IN(12) => B_ID2EXE_12_port, PAD_IN(11) => 
                           B_ID2EXE_11_port, PAD_IN(10) => B_ID2EXE_10_port, 
                           PAD_IN(9) => B_ID2EXE_9_port, PAD_IN(8) => 
                           B_ID2EXE_8_port, PAD_IN(7) => B_ID2EXE_7_port, 
                           PAD_IN(6) => B_ID2EXE_6_port, PAD_IN(5) => 
                           B_ID2EXE_5_port, PAD_IN(4) => B_ID2EXE_4_port, 
                           PAD_IN(3) => B_ID2EXE_3_port, PAD_IN(2) => 
                           B_ID2EXE_2_port, PAD_IN(1) => B_ID2EXE_1_port, 
                           PAD_IN(0) => B_ID2EXE_0_port, IR2_IN(4) => 
                           IR_ID2EXE_4_port, IR2_IN(3) => IR_ID2EXE_3_port, 
                           IR2_IN(2) => IR_ID2EXE_2_port, IR2_IN(1) => 
                           IR_ID2EXE_1_port, IR2_IN(0) => IR_ID2EXE_0_port, 
                           NPC2_OUT(31) => NPC_EXE2MEM_31_port, NPC2_OUT(30) =>
                           NPC_EXE2MEM_30_port, NPC2_OUT(29) => 
                           NPC_EXE2MEM_29_port, NPC2_OUT(28) => 
                           NPC_EXE2MEM_28_port, NPC2_OUT(27) => 
                           NPC_EXE2MEM_27_port, NPC2_OUT(26) => 
                           NPC_EXE2MEM_26_port, NPC2_OUT(25) => 
                           NPC_EXE2MEM_25_port, NPC2_OUT(24) => 
                           NPC_EXE2MEM_24_port, NPC2_OUT(23) => 
                           NPC_EXE2MEM_23_port, NPC2_OUT(22) => 
                           NPC_EXE2MEM_22_port, NPC2_OUT(21) => 
                           NPC_EXE2MEM_21_port, NPC2_OUT(20) => 
                           NPC_EXE2MEM_20_port, NPC2_OUT(19) => 
                           NPC_EXE2MEM_19_port, NPC2_OUT(18) => 
                           NPC_EXE2MEM_18_port, NPC2_OUT(17) => 
                           NPC_EXE2MEM_17_port, NPC2_OUT(16) => 
                           NPC_EXE2MEM_16_port, NPC2_OUT(15) => 
                           NPC_EXE2MEM_15_port, NPC2_OUT(14) => 
                           NPC_EXE2MEM_14_port, NPC2_OUT(13) => 
                           NPC_EXE2MEM_13_port, NPC2_OUT(12) => 
                           NPC_EXE2MEM_12_port, NPC2_OUT(11) => 
                           NPC_EXE2MEM_11_port, NPC2_OUT(10) => 
                           NPC_EXE2MEM_10_port, NPC2_OUT(9) => 
                           NPC_EXE2MEM_9_port, NPC2_OUT(8) => 
                           NPC_EXE2MEM_8_port, NPC2_OUT(7) => 
                           NPC_EXE2MEM_7_port, NPC2_OUT(6) => 
                           NPC_EXE2MEM_6_port, NPC2_OUT(5) => 
                           NPC_EXE2MEM_5_port, NPC2_OUT(4) => 
                           NPC_EXE2MEM_4_port, NPC2_OUT(3) => 
                           NPC_EXE2MEM_3_port, NPC2_OUT(2) => 
                           NPC_EXE2MEM_2_port, NPC2_OUT(1) => 
                           NPC_EXE2MEM_1_port, NPC2_OUT(0) => 
                           NPC_EXE2MEM_0_port, ZERO_OP_OUT => ZOP_EXE2MEM, 
                           ALU_OUT(31) => ALU_EXE2MEM_31_port, ALU_OUT(30) => 
                           ALU_EXE2MEM_30_port, ALU_OUT(29) => 
                           ALU_EXE2MEM_29_port, ALU_OUT(28) => 
                           ALU_EXE2MEM_28_port, ALU_OUT(27) => 
                           ALU_EXE2MEM_27_port, ALU_OUT(26) => 
                           ALU_EXE2MEM_26_port, ALU_OUT(25) => 
                           ALU_EXE2MEM_25_port, ALU_OUT(24) => 
                           ALU_EXE2MEM_24_port, ALU_OUT(23) => 
                           ALU_EXE2MEM_23_port, ALU_OUT(22) => 
                           ALU_EXE2MEM_22_port, ALU_OUT(21) => 
                           ALU_EXE2MEM_21_port, ALU_OUT(20) => 
                           ALU_EXE2MEM_20_port, ALU_OUT(19) => 
                           ALU_EXE2MEM_19_port, ALU_OUT(18) => 
                           ALU_EXE2MEM_18_port, ALU_OUT(17) => 
                           ALU_EXE2MEM_17_port, ALU_OUT(16) => 
                           ALU_EXE2MEM_16_port, ALU_OUT(15) => 
                           ALU_EXE2MEM_15_port, ALU_OUT(14) => 
                           ALU_EXE2MEM_14_port, ALU_OUT(13) => 
                           ALU_EXE2MEM_13_port, ALU_OUT(12) => 
                           ALU_EXE2MEM_12_port, ALU_OUT(11) => 
                           ALU_EXE2MEM_11_port, ALU_OUT(10) => 
                           ALU_EXE2MEM_10_port, ALU_OUT(9) => 
                           ALU_EXE2MEM_9_port, ALU_OUT(8) => ALU_EXE2MEM_8_port
                           , ALU_OUT(7) => ALU_EXE2MEM_7_port, ALU_OUT(6) => 
                           ALU_EXE2MEM_6_port, ALU_OUT(5) => ALU_EXE2MEM_5_port
                           , ALU_OUT(4) => ALU_EXE2MEM_4_port, ALU_OUT(3) => 
                           ALU_EXE2MEM_3_port, ALU_OUT(2) => ALU_EXE2MEM_2_port
                           , ALU_OUT(1) => ALU_EXE2MEM_1_port, ALU_OUT(0) => 
                           ALU_EXE2MEM_0_port, PAD_OUT(31) => 
                           PAD_EXE2MEM_31_port, PAD_OUT(30) => 
                           PAD_EXE2MEM_30_port, PAD_OUT(29) => 
                           PAD_EXE2MEM_29_port, PAD_OUT(28) => 
                           PAD_EXE2MEM_28_port, PAD_OUT(27) => 
                           PAD_EXE2MEM_27_port, PAD_OUT(26) => 
                           PAD_EXE2MEM_26_port, PAD_OUT(25) => 
                           PAD_EXE2MEM_25_port, PAD_OUT(24) => 
                           PAD_EXE2MEM_24_port, PAD_OUT(23) => 
                           PAD_EXE2MEM_23_port, PAD_OUT(22) => 
                           PAD_EXE2MEM_22_port, PAD_OUT(21) => 
                           PAD_EXE2MEM_21_port, PAD_OUT(20) => 
                           PAD_EXE2MEM_20_port, PAD_OUT(19) => 
                           PAD_EXE2MEM_19_port, PAD_OUT(18) => 
                           PAD_EXE2MEM_18_port, PAD_OUT(17) => 
                           PAD_EXE2MEM_17_port, PAD_OUT(16) => 
                           PAD_EXE2MEM_16_port, PAD_OUT(15) => 
                           PAD_EXE2MEM_15_port, PAD_OUT(14) => 
                           PAD_EXE2MEM_14_port, PAD_OUT(13) => 
                           PAD_EXE2MEM_13_port, PAD_OUT(12) => 
                           PAD_EXE2MEM_12_port, PAD_OUT(11) => 
                           PAD_EXE2MEM_11_port, PAD_OUT(10) => 
                           PAD_EXE2MEM_10_port, PAD_OUT(9) => 
                           PAD_EXE2MEM_9_port, PAD_OUT(8) => PAD_EXE2MEM_8_port
                           , PAD_OUT(7) => PAD_EXE2MEM_7_port, PAD_OUT(6) => 
                           PAD_EXE2MEM_6_port, PAD_OUT(5) => PAD_EXE2MEM_5_port
                           , PAD_OUT(4) => PAD_EXE2MEM_4_port, PAD_OUT(3) => 
                           PAD_EXE2MEM_3_port, PAD_OUT(2) => PAD_EXE2MEM_2_port
                           , PAD_OUT(1) => PAD_EXE2MEM_1_port, PAD_OUT(0) => 
                           PAD_EXE2MEM_0_port, IR2_OUT(4) => IR_EXE2MEM_4_port,
                           IR2_OUT(3) => IR_EXE2MEM_3_port, IR2_OUT(2) => 
                           IR_EXE2MEM_2_port, IR2_OUT(1) => IR_EXE2MEM_1_port, 
                           IR2_OUT(0) => IR_EXE2MEM_0_port, N_FLAG => n_2208, 
                           Z_FLAG => n_2209, C_FLAG => n_2210, V_FLAG => n_2211
                           );
   MEMORY : MEM_STAGE_N_BITS_DATA32_RF_ADDR5 port map( CLK => CLK, RST => RST, 
                           MEM_OUTREG_EN => MEM_OUTREG_EN, ZERO_PADDING4 => 
                           ZERO_PADDING4, MEM_OUT_SEL => MEM_OUT_SEL, 
                           BYTE_LEN_IN(1) => BYTE_LEN_IN(1), BYTE_LEN_IN(0) => 
                           BYTE_LEN_IN(0), DRAM_WE => DRAM_WE, DRAM_WE_OUT => 
                           DRAM_WE_OUT, BYTE_LEN_OUT(1) => BYTE_LEN_OUT(1), 
                           BYTE_LEN_OUT(0) => BYTE_LEN_OUT(0), BRA_IN => 
                           ZOP_EXE2MEM, JUMP_MUX_IN_0(31) => 
                           NPC_IF2ID_MEM_31_port, JUMP_MUX_IN_0(30) => 
                           NPC_IF2ID_MEM_30_port, JUMP_MUX_IN_0(29) => 
                           NPC_IF2ID_MEM_29_port, JUMP_MUX_IN_0(28) => 
                           NPC_IF2ID_MEM_28_port, JUMP_MUX_IN_0(27) => 
                           NPC_IF2ID_MEM_27_port, JUMP_MUX_IN_0(26) => 
                           NPC_IF2ID_MEM_26_port, JUMP_MUX_IN_0(25) => 
                           NPC_IF2ID_MEM_25_port, JUMP_MUX_IN_0(24) => 
                           NPC_IF2ID_MEM_24_port, JUMP_MUX_IN_0(23) => 
                           NPC_IF2ID_MEM_23_port, JUMP_MUX_IN_0(22) => 
                           NPC_IF2ID_MEM_22_port, JUMP_MUX_IN_0(21) => 
                           NPC_IF2ID_MEM_21_port, JUMP_MUX_IN_0(20) => 
                           NPC_IF2ID_MEM_20_port, JUMP_MUX_IN_0(19) => 
                           NPC_IF2ID_MEM_19_port, JUMP_MUX_IN_0(18) => 
                           NPC_IF2ID_MEM_18_port, JUMP_MUX_IN_0(17) => 
                           NPC_IF2ID_MEM_17_port, JUMP_MUX_IN_0(16) => 
                           NPC_IF2ID_MEM_16_port, JUMP_MUX_IN_0(15) => 
                           NPC_IF2ID_MEM_15_port, JUMP_MUX_IN_0(14) => 
                           NPC_IF2ID_MEM_14_port, JUMP_MUX_IN_0(13) => 
                           NPC_IF2ID_MEM_13_port, JUMP_MUX_IN_0(12) => 
                           NPC_IF2ID_MEM_12_port, JUMP_MUX_IN_0(11) => 
                           NPC_IF2ID_MEM_11_port, JUMP_MUX_IN_0(10) => 
                           NPC_IF2ID_MEM_10_port, JUMP_MUX_IN_0(9) => 
                           NPC_IF2ID_MEM_9_port, JUMP_MUX_IN_0(8) => 
                           NPC_IF2ID_MEM_8_port, JUMP_MUX_IN_0(7) => 
                           NPC_IF2ID_MEM_7_port, JUMP_MUX_IN_0(6) => 
                           NPC_IF2ID_MEM_6_port, JUMP_MUX_IN_0(5) => 
                           NPC_IF2ID_MEM_5_port, JUMP_MUX_IN_0(4) => 
                           NPC_IF2ID_MEM_4_port, JUMP_MUX_IN_0(3) => 
                           NPC_IF2ID_MEM_3_port, JUMP_MUX_IN_0(2) => 
                           NPC_IF2ID_MEM_2_port, JUMP_MUX_IN_0(1) => 
                           NPC_IF2ID_MEM_1_port, JUMP_MUX_IN_0(0) => 
                           NPC_IF2ID_MEM_0_port, ALU_OUTPUT_IN(31) => 
                           ALU_EXE2MEM_31_port, ALU_OUTPUT_IN(30) => 
                           ALU_EXE2MEM_30_port, ALU_OUTPUT_IN(29) => 
                           ALU_EXE2MEM_29_port, ALU_OUTPUT_IN(28) => 
                           ALU_EXE2MEM_28_port, ALU_OUTPUT_IN(27) => 
                           ALU_EXE2MEM_27_port, ALU_OUTPUT_IN(26) => 
                           ALU_EXE2MEM_26_port, ALU_OUTPUT_IN(25) => 
                           ALU_EXE2MEM_25_port, ALU_OUTPUT_IN(24) => 
                           ALU_EXE2MEM_24_port, ALU_OUTPUT_IN(23) => 
                           ALU_EXE2MEM_23_port, ALU_OUTPUT_IN(22) => 
                           ALU_EXE2MEM_22_port, ALU_OUTPUT_IN(21) => 
                           ALU_EXE2MEM_21_port, ALU_OUTPUT_IN(20) => 
                           ALU_EXE2MEM_20_port, ALU_OUTPUT_IN(19) => 
                           ALU_EXE2MEM_19_port, ALU_OUTPUT_IN(18) => 
                           ALU_EXE2MEM_18_port, ALU_OUTPUT_IN(17) => 
                           ALU_EXE2MEM_17_port, ALU_OUTPUT_IN(16) => 
                           ALU_EXE2MEM_16_port, ALU_OUTPUT_IN(15) => 
                           ALU_EXE2MEM_15_port, ALU_OUTPUT_IN(14) => 
                           ALU_EXE2MEM_14_port, ALU_OUTPUT_IN(13) => 
                           ALU_EXE2MEM_13_port, ALU_OUTPUT_IN(12) => 
                           ALU_EXE2MEM_12_port, ALU_OUTPUT_IN(11) => 
                           ALU_EXE2MEM_11_port, ALU_OUTPUT_IN(10) => 
                           ALU_EXE2MEM_10_port, ALU_OUTPUT_IN(9) => 
                           ALU_EXE2MEM_9_port, ALU_OUTPUT_IN(8) => 
                           ALU_EXE2MEM_8_port, ALU_OUTPUT_IN(7) => 
                           ALU_EXE2MEM_7_port, ALU_OUTPUT_IN(6) => 
                           ALU_EXE2MEM_6_port, ALU_OUTPUT_IN(5) => 
                           ALU_EXE2MEM_5_port, ALU_OUTPUT_IN(4) => 
                           ALU_EXE2MEM_4_port, ALU_OUTPUT_IN(3) => 
                           ALU_EXE2MEM_3_port, ALU_OUTPUT_IN(2) => 
                           ALU_EXE2MEM_2_port, ALU_OUTPUT_IN(1) => 
                           ALU_EXE2MEM_1_port, ALU_OUTPUT_IN(0) => 
                           ALU_EXE2MEM_0_port, MEM_DATA_IN(31) => 
                           PAD_EXE2MEM_31_port, MEM_DATA_IN(30) => 
                           PAD_EXE2MEM_30_port, MEM_DATA_IN(29) => 
                           PAD_EXE2MEM_29_port, MEM_DATA_IN(28) => 
                           PAD_EXE2MEM_28_port, MEM_DATA_IN(27) => 
                           PAD_EXE2MEM_27_port, MEM_DATA_IN(26) => 
                           PAD_EXE2MEM_26_port, MEM_DATA_IN(25) => 
                           PAD_EXE2MEM_25_port, MEM_DATA_IN(24) => 
                           PAD_EXE2MEM_24_port, MEM_DATA_IN(23) => 
                           PAD_EXE2MEM_23_port, MEM_DATA_IN(22) => 
                           PAD_EXE2MEM_22_port, MEM_DATA_IN(21) => 
                           PAD_EXE2MEM_21_port, MEM_DATA_IN(20) => 
                           PAD_EXE2MEM_20_port, MEM_DATA_IN(19) => 
                           PAD_EXE2MEM_19_port, MEM_DATA_IN(18) => 
                           PAD_EXE2MEM_18_port, MEM_DATA_IN(17) => 
                           PAD_EXE2MEM_17_port, MEM_DATA_IN(16) => 
                           PAD_EXE2MEM_16_port, MEM_DATA_IN(15) => 
                           PAD_EXE2MEM_15_port, MEM_DATA_IN(14) => 
                           PAD_EXE2MEM_14_port, MEM_DATA_IN(13) => 
                           PAD_EXE2MEM_13_port, MEM_DATA_IN(12) => 
                           PAD_EXE2MEM_12_port, MEM_DATA_IN(11) => 
                           PAD_EXE2MEM_11_port, MEM_DATA_IN(10) => 
                           PAD_EXE2MEM_10_port, MEM_DATA_IN(9) => 
                           PAD_EXE2MEM_9_port, MEM_DATA_IN(8) => 
                           PAD_EXE2MEM_8_port, MEM_DATA_IN(7) => 
                           PAD_EXE2MEM_7_port, MEM_DATA_IN(6) => 
                           PAD_EXE2MEM_6_port, MEM_DATA_IN(5) => 
                           PAD_EXE2MEM_5_port, MEM_DATA_IN(4) => 
                           PAD_EXE2MEM_4_port, MEM_DATA_IN(3) => 
                           PAD_EXE2MEM_3_port, MEM_DATA_IN(2) => 
                           PAD_EXE2MEM_2_port, MEM_DATA_IN(1) => 
                           PAD_EXE2MEM_1_port, MEM_DATA_IN(0) => 
                           PAD_EXE2MEM_0_port, MEM_DATA_OUT_INT(31) => 
                           MEM_DATA_OUT_INT(31), MEM_DATA_OUT_INT(30) => 
                           MEM_DATA_OUT_INT(30), MEM_DATA_OUT_INT(29) => 
                           MEM_DATA_OUT_INT(29), MEM_DATA_OUT_INT(28) => 
                           MEM_DATA_OUT_INT(28), MEM_DATA_OUT_INT(27) => 
                           MEM_DATA_OUT_INT(27), MEM_DATA_OUT_INT(26) => 
                           MEM_DATA_OUT_INT(26), MEM_DATA_OUT_INT(25) => 
                           MEM_DATA_OUT_INT(25), MEM_DATA_OUT_INT(24) => 
                           MEM_DATA_OUT_INT(24), MEM_DATA_OUT_INT(23) => 
                           MEM_DATA_OUT_INT(23), MEM_DATA_OUT_INT(22) => 
                           MEM_DATA_OUT_INT(22), MEM_DATA_OUT_INT(21) => 
                           MEM_DATA_OUT_INT(21), MEM_DATA_OUT_INT(20) => 
                           MEM_DATA_OUT_INT(20), MEM_DATA_OUT_INT(19) => 
                           MEM_DATA_OUT_INT(19), MEM_DATA_OUT_INT(18) => 
                           MEM_DATA_OUT_INT(18), MEM_DATA_OUT_INT(17) => 
                           MEM_DATA_OUT_INT(17), MEM_DATA_OUT_INT(16) => 
                           MEM_DATA_OUT_INT(16), MEM_DATA_OUT_INT(15) => 
                           MEM_DATA_OUT_INT(15), MEM_DATA_OUT_INT(14) => 
                           MEM_DATA_OUT_INT(14), MEM_DATA_OUT_INT(13) => 
                           MEM_DATA_OUT_INT(13), MEM_DATA_OUT_INT(12) => 
                           MEM_DATA_OUT_INT(12), MEM_DATA_OUT_INT(11) => 
                           MEM_DATA_OUT_INT(11), MEM_DATA_OUT_INT(10) => 
                           MEM_DATA_OUT_INT(10), MEM_DATA_OUT_INT(9) => 
                           MEM_DATA_OUT_INT(9), MEM_DATA_OUT_INT(8) => 
                           MEM_DATA_OUT_INT(8), MEM_DATA_OUT_INT(7) => 
                           MEM_DATA_OUT_INT(7), MEM_DATA_OUT_INT(6) => 
                           MEM_DATA_OUT_INT(6), MEM_DATA_OUT_INT(5) => 
                           MEM_DATA_OUT_INT(5), MEM_DATA_OUT_INT(4) => 
                           MEM_DATA_OUT_INT(4), MEM_DATA_OUT_INT(3) => 
                           MEM_DATA_OUT_INT(3), MEM_DATA_OUT_INT(2) => 
                           MEM_DATA_OUT_INT(2), MEM_DATA_OUT_INT(1) => 
                           MEM_DATA_OUT_INT(1), MEM_DATA_OUT_INT(0) => 
                           MEM_DATA_OUT_INT(0), NPC_IN(31) => 
                           NPC_EXE2MEM_31_port, NPC_IN(30) => 
                           NPC_EXE2MEM_30_port, NPC_IN(29) => 
                           NPC_EXE2MEM_29_port, NPC_IN(28) => 
                           NPC_EXE2MEM_28_port, NPC_IN(27) => 
                           NPC_EXE2MEM_27_port, NPC_IN(26) => 
                           NPC_EXE2MEM_26_port, NPC_IN(25) => 
                           NPC_EXE2MEM_25_port, NPC_IN(24) => 
                           NPC_EXE2MEM_24_port, NPC_IN(23) => 
                           NPC_EXE2MEM_23_port, NPC_IN(22) => 
                           NPC_EXE2MEM_22_port, NPC_IN(21) => 
                           NPC_EXE2MEM_21_port, NPC_IN(20) => 
                           NPC_EXE2MEM_20_port, NPC_IN(19) => 
                           NPC_EXE2MEM_19_port, NPC_IN(18) => 
                           NPC_EXE2MEM_18_port, NPC_IN(17) => 
                           NPC_EXE2MEM_17_port, NPC_IN(16) => 
                           NPC_EXE2MEM_16_port, NPC_IN(15) => 
                           NPC_EXE2MEM_15_port, NPC_IN(14) => 
                           NPC_EXE2MEM_14_port, NPC_IN(13) => 
                           NPC_EXE2MEM_13_port, NPC_IN(12) => 
                           NPC_EXE2MEM_12_port, NPC_IN(11) => 
                           NPC_EXE2MEM_11_port, NPC_IN(10) => 
                           NPC_EXE2MEM_10_port, NPC_IN(9) => NPC_EXE2MEM_9_port
                           , NPC_IN(8) => NPC_EXE2MEM_8_port, NPC_IN(7) => 
                           NPC_EXE2MEM_7_port, NPC_IN(6) => NPC_EXE2MEM_6_port,
                           NPC_IN(5) => NPC_EXE2MEM_5_port, NPC_IN(4) => 
                           NPC_EXE2MEM_4_port, NPC_IN(3) => NPC_EXE2MEM_3_port,
                           NPC_IN(2) => NPC_EXE2MEM_2_port, NPC_IN(1) => 
                           NPC_EXE2MEM_1_port, NPC_IN(0) => NPC_EXE2MEM_0_port,
                           IR_IN(4) => IR_EXE2MEM_4_port, IR_IN(3) => 
                           IR_EXE2MEM_3_port, IR_IN(2) => IR_EXE2MEM_2_port, 
                           IR_IN(1) => IR_EXE2MEM_1_port, IR_IN(0) => 
                           IR_EXE2MEM_0_port, IR_OUT(4) => IR_MEM2WB_4_port, 
                           IR_OUT(3) => IR_MEM2WB_3_port, IR_OUT(2) => 
                           IR_MEM2WB_2_port, IR_OUT(1) => IR_MEM2WB_1_port, 
                           IR_OUT(0) => IR_MEM2WB_0_port, NPC_OUT(31) => 
                           NPC_MEM2WB_31_port, NPC_OUT(30) => 
                           NPC_MEM2WB_30_port, NPC_OUT(29) => 
                           NPC_MEM2WB_29_port, NPC_OUT(28) => 
                           NPC_MEM2WB_28_port, NPC_OUT(27) => 
                           NPC_MEM2WB_27_port, NPC_OUT(26) => 
                           NPC_MEM2WB_26_port, NPC_OUT(25) => 
                           NPC_MEM2WB_25_port, NPC_OUT(24) => 
                           NPC_MEM2WB_24_port, NPC_OUT(23) => 
                           NPC_MEM2WB_23_port, NPC_OUT(22) => 
                           NPC_MEM2WB_22_port, NPC_OUT(21) => 
                           NPC_MEM2WB_21_port, NPC_OUT(20) => 
                           NPC_MEM2WB_20_port, NPC_OUT(19) => 
                           NPC_MEM2WB_19_port, NPC_OUT(18) => 
                           NPC_MEM2WB_18_port, NPC_OUT(17) => 
                           NPC_MEM2WB_17_port, NPC_OUT(16) => 
                           NPC_MEM2WB_16_port, NPC_OUT(15) => 
                           NPC_MEM2WB_15_port, NPC_OUT(14) => 
                           NPC_MEM2WB_14_port, NPC_OUT(13) => 
                           NPC_MEM2WB_13_port, NPC_OUT(12) => 
                           NPC_MEM2WB_12_port, NPC_OUT(11) => 
                           NPC_MEM2WB_11_port, NPC_OUT(10) => 
                           NPC_MEM2WB_10_port, NPC_OUT(9) => NPC_MEM2WB_9_port,
                           NPC_OUT(8) => NPC_MEM2WB_8_port, NPC_OUT(7) => 
                           NPC_MEM2WB_7_port, NPC_OUT(6) => NPC_MEM2WB_6_port, 
                           NPC_OUT(5) => NPC_MEM2WB_5_port, NPC_OUT(4) => 
                           NPC_MEM2WB_4_port, NPC_OUT(3) => NPC_MEM2WB_3_port, 
                           NPC_OUT(2) => NPC_MEM2WB_2_port, NPC_OUT(1) => 
                           NPC_MEM2WB_1_port, NPC_OUT(0) => NPC_MEM2WB_0_port, 
                           MEM_ADDR_OUT(31) => MEM_ADDR_OUT(31), 
                           MEM_ADDR_OUT(30) => MEM_ADDR_OUT(30), 
                           MEM_ADDR_OUT(29) => MEM_ADDR_OUT(29), 
                           MEM_ADDR_OUT(28) => MEM_ADDR_OUT(28), 
                           MEM_ADDR_OUT(27) => MEM_ADDR_OUT(27), 
                           MEM_ADDR_OUT(26) => MEM_ADDR_OUT(26), 
                           MEM_ADDR_OUT(25) => MEM_ADDR_OUT(25), 
                           MEM_ADDR_OUT(24) => MEM_ADDR_OUT(24), 
                           MEM_ADDR_OUT(23) => MEM_ADDR_OUT(23), 
                           MEM_ADDR_OUT(22) => MEM_ADDR_OUT(22), 
                           MEM_ADDR_OUT(21) => MEM_ADDR_OUT(21), 
                           MEM_ADDR_OUT(20) => MEM_ADDR_OUT(20), 
                           MEM_ADDR_OUT(19) => MEM_ADDR_OUT(19), 
                           MEM_ADDR_OUT(18) => MEM_ADDR_OUT(18), 
                           MEM_ADDR_OUT(17) => MEM_ADDR_OUT(17), 
                           MEM_ADDR_OUT(16) => MEM_ADDR_OUT(16), 
                           MEM_ADDR_OUT(15) => MEM_ADDR_OUT(15), 
                           MEM_ADDR_OUT(14) => MEM_ADDR_OUT(14), 
                           MEM_ADDR_OUT(13) => MEM_ADDR_OUT(13), 
                           MEM_ADDR_OUT(12) => MEM_ADDR_OUT(12), 
                           MEM_ADDR_OUT(11) => MEM_ADDR_OUT(11), 
                           MEM_ADDR_OUT(10) => MEM_ADDR_OUT(10), 
                           MEM_ADDR_OUT(9) => MEM_ADDR_OUT(9), MEM_ADDR_OUT(8) 
                           => MEM_ADDR_OUT(8), MEM_ADDR_OUT(7) => 
                           MEM_ADDR_OUT(7), MEM_ADDR_OUT(6) => MEM_ADDR_OUT(6),
                           MEM_ADDR_OUT(5) => MEM_ADDR_OUT(5), MEM_ADDR_OUT(4) 
                           => MEM_ADDR_OUT(4), MEM_ADDR_OUT(3) => 
                           MEM_ADDR_OUT(3), MEM_ADDR_OUT(2) => MEM_ADDR_OUT(2),
                           MEM_ADDR_OUT(1) => MEM_ADDR_OUT(1), MEM_ADDR_OUT(0) 
                           => MEM_ADDR_OUT(0), MEM_DATA_IN_PRIME(31) => 
                           MEM_DATA_IN_PRIME(31), MEM_DATA_IN_PRIME(30) => 
                           MEM_DATA_IN_PRIME(30), MEM_DATA_IN_PRIME(29) => 
                           MEM_DATA_IN_PRIME(29), MEM_DATA_IN_PRIME(28) => 
                           MEM_DATA_IN_PRIME(28), MEM_DATA_IN_PRIME(27) => 
                           MEM_DATA_IN_PRIME(27), MEM_DATA_IN_PRIME(26) => 
                           MEM_DATA_IN_PRIME(26), MEM_DATA_IN_PRIME(25) => 
                           MEM_DATA_IN_PRIME(25), MEM_DATA_IN_PRIME(24) => 
                           MEM_DATA_IN_PRIME(24), MEM_DATA_IN_PRIME(23) => 
                           MEM_DATA_IN_PRIME(23), MEM_DATA_IN_PRIME(22) => 
                           MEM_DATA_IN_PRIME(22), MEM_DATA_IN_PRIME(21) => 
                           MEM_DATA_IN_PRIME(21), MEM_DATA_IN_PRIME(20) => 
                           MEM_DATA_IN_PRIME(20), MEM_DATA_IN_PRIME(19) => 
                           MEM_DATA_IN_PRIME(19), MEM_DATA_IN_PRIME(18) => 
                           MEM_DATA_IN_PRIME(18), MEM_DATA_IN_PRIME(17) => 
                           MEM_DATA_IN_PRIME(17), MEM_DATA_IN_PRIME(16) => 
                           MEM_DATA_IN_PRIME(16), MEM_DATA_IN_PRIME(15) => 
                           MEM_DATA_IN_PRIME(15), MEM_DATA_IN_PRIME(14) => 
                           MEM_DATA_IN_PRIME(14), MEM_DATA_IN_PRIME(13) => 
                           MEM_DATA_IN_PRIME(13), MEM_DATA_IN_PRIME(12) => 
                           MEM_DATA_IN_PRIME(12), MEM_DATA_IN_PRIME(11) => 
                           MEM_DATA_IN_PRIME(11), MEM_DATA_IN_PRIME(10) => 
                           MEM_DATA_IN_PRIME(10), MEM_DATA_IN_PRIME(9) => 
                           MEM_DATA_IN_PRIME(9), MEM_DATA_IN_PRIME(8) => 
                           MEM_DATA_IN_PRIME(8), MEM_DATA_IN_PRIME(7) => 
                           MEM_DATA_IN_PRIME(7), MEM_DATA_IN_PRIME(6) => 
                           MEM_DATA_IN_PRIME(6), MEM_DATA_IN_PRIME(5) => 
                           MEM_DATA_IN_PRIME(5), MEM_DATA_IN_PRIME(4) => 
                           MEM_DATA_IN_PRIME(4), MEM_DATA_IN_PRIME(3) => 
                           MEM_DATA_IN_PRIME(3), MEM_DATA_IN_PRIME(2) => 
                           MEM_DATA_IN_PRIME(2), MEM_DATA_IN_PRIME(1) => 
                           MEM_DATA_IN_PRIME(1), MEM_DATA_IN_PRIME(0) => 
                           MEM_DATA_IN_PRIME(0), ALU_OUTPUT_OUT(31) => 
                           ALU_MEM2WB_31_port, ALU_OUTPUT_OUT(30) => 
                           ALU_MEM2WB_30_port, ALU_OUTPUT_OUT(29) => 
                           ALU_MEM2WB_29_port, ALU_OUTPUT_OUT(28) => 
                           ALU_MEM2WB_28_port, ALU_OUTPUT_OUT(27) => 
                           ALU_MEM2WB_27_port, ALU_OUTPUT_OUT(26) => 
                           ALU_MEM2WB_26_port, ALU_OUTPUT_OUT(25) => 
                           ALU_MEM2WB_25_port, ALU_OUTPUT_OUT(24) => 
                           ALU_MEM2WB_24_port, ALU_OUTPUT_OUT(23) => 
                           ALU_MEM2WB_23_port, ALU_OUTPUT_OUT(22) => 
                           ALU_MEM2WB_22_port, ALU_OUTPUT_OUT(21) => 
                           ALU_MEM2WB_21_port, ALU_OUTPUT_OUT(20) => 
                           ALU_MEM2WB_20_port, ALU_OUTPUT_OUT(19) => 
                           ALU_MEM2WB_19_port, ALU_OUTPUT_OUT(18) => 
                           ALU_MEM2WB_18_port, ALU_OUTPUT_OUT(17) => 
                           ALU_MEM2WB_17_port, ALU_OUTPUT_OUT(16) => 
                           ALU_MEM2WB_16_port, ALU_OUTPUT_OUT(15) => 
                           ALU_MEM2WB_15_port, ALU_OUTPUT_OUT(14) => 
                           ALU_MEM2WB_14_port, ALU_OUTPUT_OUT(13) => 
                           ALU_MEM2WB_13_port, ALU_OUTPUT_OUT(12) => 
                           ALU_MEM2WB_12_port, ALU_OUTPUT_OUT(11) => 
                           ALU_MEM2WB_11_port, ALU_OUTPUT_OUT(10) => 
                           ALU_MEM2WB_10_port, ALU_OUTPUT_OUT(9) => 
                           ALU_MEM2WB_9_port, ALU_OUTPUT_OUT(8) => 
                           ALU_MEM2WB_8_port, ALU_OUTPUT_OUT(7) => 
                           ALU_MEM2WB_7_port, ALU_OUTPUT_OUT(6) => 
                           ALU_MEM2WB_6_port, ALU_OUTPUT_OUT(5) => 
                           ALU_MEM2WB_5_port, ALU_OUTPUT_OUT(4) => 
                           ALU_MEM2WB_4_port, ALU_OUTPUT_OUT(3) => 
                           ALU_MEM2WB_3_port, ALU_OUTPUT_OUT(2) => 
                           ALU_MEM2WB_2_port, ALU_OUTPUT_OUT(1) => 
                           ALU_MEM2WB_1_port, ALU_OUTPUT_OUT(0) => 
                           ALU_MEM2WB_0_port, MEM_DATA_OUT(31) => 
                           MEM_MEM2WB_31_port, MEM_DATA_OUT(30) => 
                           MEM_MEM2WB_30_port, MEM_DATA_OUT(29) => 
                           MEM_MEM2WB_29_port, MEM_DATA_OUT(28) => 
                           MEM_MEM2WB_28_port, MEM_DATA_OUT(27) => 
                           MEM_MEM2WB_27_port, MEM_DATA_OUT(26) => 
                           MEM_MEM2WB_26_port, MEM_DATA_OUT(25) => 
                           MEM_MEM2WB_25_port, MEM_DATA_OUT(24) => 
                           MEM_MEM2WB_24_port, MEM_DATA_OUT(23) => 
                           MEM_MEM2WB_23_port, MEM_DATA_OUT(22) => 
                           MEM_MEM2WB_22_port, MEM_DATA_OUT(21) => 
                           MEM_MEM2WB_21_port, MEM_DATA_OUT(20) => 
                           MEM_MEM2WB_20_port, MEM_DATA_OUT(19) => 
                           MEM_MEM2WB_19_port, MEM_DATA_OUT(18) => 
                           MEM_MEM2WB_18_port, MEM_DATA_OUT(17) => 
                           MEM_MEM2WB_17_port, MEM_DATA_OUT(16) => 
                           MEM_MEM2WB_16_port, MEM_DATA_OUT(15) => 
                           MEM_MEM2WB_15_port, MEM_DATA_OUT(14) => 
                           MEM_MEM2WB_14_port, MEM_DATA_OUT(13) => 
                           MEM_MEM2WB_13_port, MEM_DATA_OUT(12) => 
                           MEM_MEM2WB_12_port, MEM_DATA_OUT(11) => 
                           MEM_MEM2WB_11_port, MEM_DATA_OUT(10) => 
                           MEM_MEM2WB_10_port, MEM_DATA_OUT(9) => 
                           MEM_MEM2WB_9_port, MEM_DATA_OUT(8) => 
                           MEM_MEM2WB_8_port, MEM_DATA_OUT(7) => 
                           MEM_MEM2WB_7_port, MEM_DATA_OUT(6) => 
                           MEM_MEM2WB_6_port, MEM_DATA_OUT(5) => 
                           MEM_MEM2WB_5_port, MEM_DATA_OUT(4) => 
                           MEM_MEM2WB_4_port, MEM_DATA_OUT(3) => 
                           MEM_MEM2WB_3_port, MEM_DATA_OUT(2) => 
                           MEM_MEM2WB_2_port, MEM_DATA_OUT(1) => 
                           MEM_MEM2WB_1_port, MEM_DATA_OUT(0) => 
                           MEM_MEM2WB_0_port, ADDR_MUX_OUT(31) => 
                           PC_MEM2IF_31_port, ADDR_MUX_OUT(30) => 
                           PC_MEM2IF_30_port, ADDR_MUX_OUT(29) => 
                           PC_MEM2IF_29_port, ADDR_MUX_OUT(28) => 
                           PC_MEM2IF_28_port, ADDR_MUX_OUT(27) => 
                           PC_MEM2IF_27_port, ADDR_MUX_OUT(26) => 
                           PC_MEM2IF_26_port, ADDR_MUX_OUT(25) => 
                           PC_MEM2IF_25_port, ADDR_MUX_OUT(24) => 
                           PC_MEM2IF_24_port, ADDR_MUX_OUT(23) => 
                           PC_MEM2IF_23_port, ADDR_MUX_OUT(22) => 
                           PC_MEM2IF_22_port, ADDR_MUX_OUT(21) => 
                           PC_MEM2IF_21_port, ADDR_MUX_OUT(20) => 
                           PC_MEM2IF_20_port, ADDR_MUX_OUT(19) => 
                           PC_MEM2IF_19_port, ADDR_MUX_OUT(18) => 
                           PC_MEM2IF_18_port, ADDR_MUX_OUT(17) => 
                           PC_MEM2IF_17_port, ADDR_MUX_OUT(16) => 
                           PC_MEM2IF_16_port, ADDR_MUX_OUT(15) => 
                           PC_MEM2IF_15_port, ADDR_MUX_OUT(14) => 
                           PC_MEM2IF_14_port, ADDR_MUX_OUT(13) => 
                           PC_MEM2IF_13_port, ADDR_MUX_OUT(12) => 
                           PC_MEM2IF_12_port, ADDR_MUX_OUT(11) => 
                           PC_MEM2IF_11_port, ADDR_MUX_OUT(10) => 
                           PC_MEM2IF_10_port, ADDR_MUX_OUT(9) => 
                           PC_MEM2IF_9_port, ADDR_MUX_OUT(8) => 
                           PC_MEM2IF_8_port, ADDR_MUX_OUT(7) => 
                           PC_MEM2IF_7_port, ADDR_MUX_OUT(6) => 
                           PC_MEM2IF_6_port, ADDR_MUX_OUT(5) => 
                           PC_MEM2IF_5_port, ADDR_MUX_OUT(4) => 
                           PC_MEM2IF_4_port, ADDR_MUX_OUT(3) => 
                           PC_MEM2IF_3_port, ADDR_MUX_OUT(2) => 
                           PC_MEM2IF_2_port, ADDR_MUX_OUT(1) => 
                           PC_MEM2IF_1_port, ADDR_MUX_OUT(0) => 
                           PC_MEM2IF_0_port);
   WRITE_BACK : WB_STAGE_N_BITS_DATA32_RF_ADDR5 port map( CLK => CLK, RST => 
                           RST, WB_LATCH_EN => WB_LATCH_EN, JAL_MUX_SEL => 
                           JAL_MUX_SEL, WB_MUX_SEL => WB_MUX_SEL, IR_IN(4) => 
                           IR_MEM2WB_4_port, IR_IN(3) => IR_MEM2WB_3_port, 
                           IR_IN(2) => IR_MEM2WB_2_port, IR_IN(1) => 
                           IR_MEM2WB_1_port, IR_IN(0) => IR_MEM2WB_0_port, 
                           MUX_IN2(31) => NPC_MEM2WB_31_port, MUX_IN2(30) => 
                           NPC_MEM2WB_30_port, MUX_IN2(29) => 
                           NPC_MEM2WB_29_port, MUX_IN2(28) => 
                           NPC_MEM2WB_28_port, MUX_IN2(27) => 
                           NPC_MEM2WB_27_port, MUX_IN2(26) => 
                           NPC_MEM2WB_26_port, MUX_IN2(25) => 
                           NPC_MEM2WB_25_port, MUX_IN2(24) => 
                           NPC_MEM2WB_24_port, MUX_IN2(23) => 
                           NPC_MEM2WB_23_port, MUX_IN2(22) => 
                           NPC_MEM2WB_22_port, MUX_IN2(21) => 
                           NPC_MEM2WB_21_port, MUX_IN2(20) => 
                           NPC_MEM2WB_20_port, MUX_IN2(19) => 
                           NPC_MEM2WB_19_port, MUX_IN2(18) => 
                           NPC_MEM2WB_18_port, MUX_IN2(17) => 
                           NPC_MEM2WB_17_port, MUX_IN2(16) => 
                           NPC_MEM2WB_16_port, MUX_IN2(15) => 
                           NPC_MEM2WB_15_port, MUX_IN2(14) => 
                           NPC_MEM2WB_14_port, MUX_IN2(13) => 
                           NPC_MEM2WB_13_port, MUX_IN2(12) => 
                           NPC_MEM2WB_12_port, MUX_IN2(11) => 
                           NPC_MEM2WB_11_port, MUX_IN2(10) => 
                           NPC_MEM2WB_10_port, MUX_IN2(9) => NPC_MEM2WB_9_port,
                           MUX_IN2(8) => NPC_MEM2WB_8_port, MUX_IN2(7) => 
                           NPC_MEM2WB_7_port, MUX_IN2(6) => NPC_MEM2WB_6_port, 
                           MUX_IN2(5) => NPC_MEM2WB_5_port, MUX_IN2(4) => 
                           NPC_MEM2WB_4_port, MUX_IN2(3) => NPC_MEM2WB_3_port, 
                           MUX_IN2(2) => NPC_MEM2WB_2_port, MUX_IN2(1) => 
                           NPC_MEM2WB_1_port, MUX_IN2(0) => NPC_MEM2WB_0_port, 
                           MUX_IN1(31) => MEM_MEM2WB_31_port, MUX_IN1(30) => 
                           MEM_MEM2WB_30_port, MUX_IN1(29) => 
                           MEM_MEM2WB_29_port, MUX_IN1(28) => 
                           MEM_MEM2WB_28_port, MUX_IN1(27) => 
                           MEM_MEM2WB_27_port, MUX_IN1(26) => 
                           MEM_MEM2WB_26_port, MUX_IN1(25) => 
                           MEM_MEM2WB_25_port, MUX_IN1(24) => 
                           MEM_MEM2WB_24_port, MUX_IN1(23) => 
                           MEM_MEM2WB_23_port, MUX_IN1(22) => 
                           MEM_MEM2WB_22_port, MUX_IN1(21) => 
                           MEM_MEM2WB_21_port, MUX_IN1(20) => 
                           MEM_MEM2WB_20_port, MUX_IN1(19) => 
                           MEM_MEM2WB_19_port, MUX_IN1(18) => 
                           MEM_MEM2WB_18_port, MUX_IN1(17) => 
                           MEM_MEM2WB_17_port, MUX_IN1(16) => 
                           MEM_MEM2WB_16_port, MUX_IN1(15) => 
                           MEM_MEM2WB_15_port, MUX_IN1(14) => 
                           MEM_MEM2WB_14_port, MUX_IN1(13) => 
                           MEM_MEM2WB_13_port, MUX_IN1(12) => 
                           MEM_MEM2WB_12_port, MUX_IN1(11) => 
                           MEM_MEM2WB_11_port, MUX_IN1(10) => 
                           MEM_MEM2WB_10_port, MUX_IN1(9) => MEM_MEM2WB_9_port,
                           MUX_IN1(8) => MEM_MEM2WB_8_port, MUX_IN1(7) => 
                           MEM_MEM2WB_7_port, MUX_IN1(6) => MEM_MEM2WB_6_port, 
                           MUX_IN1(5) => MEM_MEM2WB_5_port, MUX_IN1(4) => 
                           MEM_MEM2WB_4_port, MUX_IN1(3) => MEM_MEM2WB_3_port, 
                           MUX_IN1(2) => MEM_MEM2WB_2_port, MUX_IN1(1) => 
                           MEM_MEM2WB_1_port, MUX_IN1(0) => MEM_MEM2WB_0_port, 
                           MUX_IN0(31) => ALU_MEM2WB_31_port, MUX_IN0(30) => 
                           ALU_MEM2WB_30_port, MUX_IN0(29) => 
                           ALU_MEM2WB_29_port, MUX_IN0(28) => 
                           ALU_MEM2WB_28_port, MUX_IN0(27) => 
                           ALU_MEM2WB_27_port, MUX_IN0(26) => 
                           ALU_MEM2WB_26_port, MUX_IN0(25) => 
                           ALU_MEM2WB_25_port, MUX_IN0(24) => 
                           ALU_MEM2WB_24_port, MUX_IN0(23) => 
                           ALU_MEM2WB_23_port, MUX_IN0(22) => 
                           ALU_MEM2WB_22_port, MUX_IN0(21) => 
                           ALU_MEM2WB_21_port, MUX_IN0(20) => 
                           ALU_MEM2WB_20_port, MUX_IN0(19) => 
                           ALU_MEM2WB_19_port, MUX_IN0(18) => 
                           ALU_MEM2WB_18_port, MUX_IN0(17) => 
                           ALU_MEM2WB_17_port, MUX_IN0(16) => 
                           ALU_MEM2WB_16_port, MUX_IN0(15) => 
                           ALU_MEM2WB_15_port, MUX_IN0(14) => 
                           ALU_MEM2WB_14_port, MUX_IN0(13) => 
                           ALU_MEM2WB_13_port, MUX_IN0(12) => 
                           ALU_MEM2WB_12_port, MUX_IN0(11) => 
                           ALU_MEM2WB_11_port, MUX_IN0(10) => 
                           ALU_MEM2WB_10_port, MUX_IN0(9) => ALU_MEM2WB_9_port,
                           MUX_IN0(8) => ALU_MEM2WB_8_port, MUX_IN0(7) => 
                           ALU_MEM2WB_7_port, MUX_IN0(6) => ALU_MEM2WB_6_port, 
                           MUX_IN0(5) => ALU_MEM2WB_5_port, MUX_IN0(4) => 
                           ALU_MEM2WB_4_port, MUX_IN0(3) => ALU_MEM2WB_3_port, 
                           MUX_IN0(2) => ALU_MEM2WB_2_port, MUX_IN0(1) => 
                           ALU_MEM2WB_1_port, MUX_IN0(0) => ALU_MEM2WB_0_port, 
                           WRT_OUT(31) => WRT_WB2ID_31_port, WRT_OUT(30) => 
                           WRT_WB2ID_30_port, WRT_OUT(29) => WRT_WB2ID_29_port,
                           WRT_OUT(28) => WRT_WB2ID_28_port, WRT_OUT(27) => 
                           WRT_WB2ID_27_port, WRT_OUT(26) => WRT_WB2ID_26_port,
                           WRT_OUT(25) => WRT_WB2ID_25_port, WRT_OUT(24) => 
                           WRT_WB2ID_24_port, WRT_OUT(23) => WRT_WB2ID_23_port,
                           WRT_OUT(22) => WRT_WB2ID_22_port, WRT_OUT(21) => 
                           WRT_WB2ID_21_port, WRT_OUT(20) => WRT_WB2ID_20_port,
                           WRT_OUT(19) => WRT_WB2ID_19_port, WRT_OUT(18) => 
                           WRT_WB2ID_18_port, WRT_OUT(17) => WRT_WB2ID_17_port,
                           WRT_OUT(16) => WRT_WB2ID_16_port, WRT_OUT(15) => 
                           WRT_WB2ID_15_port, WRT_OUT(14) => WRT_WB2ID_14_port,
                           WRT_OUT(13) => WRT_WB2ID_13_port, WRT_OUT(12) => 
                           WRT_WB2ID_12_port, WRT_OUT(11) => WRT_WB2ID_11_port,
                           WRT_OUT(10) => WRT_WB2ID_10_port, WRT_OUT(9) => 
                           WRT_WB2ID_9_port, WRT_OUT(8) => WRT_WB2ID_8_port, 
                           WRT_OUT(7) => WRT_WB2ID_7_port, WRT_OUT(6) => 
                           WRT_WB2ID_6_port, WRT_OUT(5) => WRT_WB2ID_5_port, 
                           WRT_OUT(4) => WRT_WB2ID_4_port, WRT_OUT(3) => 
                           WRT_WB2ID_3_port, WRT_OUT(2) => WRT_WB2ID_2_port, 
                           WRT_OUT(1) => WRT_WB2ID_1_port, WRT_OUT(0) => 
                           WRT_WB2ID_0_port, IR_OUT(4) => IR_WB2ID_4_port, 
                           IR_OUT(3) => IR_WB2ID_3_port, IR_OUT(2) => 
                           IR_WB2ID_2_port, IR_OUT(1) => IR_WB2ID_1_port, 
                           IR_OUT(0) => IR_WB2ID_0_port);

end SYN_PIPELINED;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clock, ResetN : in std_logic;  Instr_In : in std_logic_vector (31 
         downto 0);  ProgCount_Out : out std_logic_vector (31 downto 0);  
         DataMem_WrEn : out std_logic;  DataMem_BLen : out std_logic_vector (1 
         downto 0);  DataMem_Addr, DataMem_Write : out std_logic_vector (31 
         downto 0);  DataMem_Read : in std_logic_vector (31 downto 0));

end DLX;

architecture SYN_PRO of DLX is

   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE22
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, 
            ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN 
            : out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 6);  
            FPU_OPCODE : out std_logic_vector (0 to 4);  PC_LATCH_EN, 
            MEM_OUTREG_EN, ZERO_PADDING4, MEM_OUT_SEL, DRAM_WE : out std_logic;
            BYTE_LEN : out std_logic_vector (1 downto 0);  WB_MUX_SEL, 
            JAL_MUX_SEL, WR_EN, WB_LATCH_EN : out std_logic);
   end component;
   
   component DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16
      port( CLK, RST, IF_LATCH_EN, PC_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, 
            RD1_EN, RD2_EN, WR_EN, ZERO_PADDING2, MUXA_SEL, MUXB_SEL, 
            EXE_OUTREG_EN, EQ_COND, JUMP_EN : in std_logic;  ALU_OPCODE : in 
            std_logic_vector (0 to 6);  MEM_OUTREG_EN, ZERO_PADDING4, 
            MEM_OUT_SEL : in std_logic;  BYTE_LEN_IN : in std_logic_vector (1 
            downto 0);  DRAM_WE : in std_logic;  DRAM_WE_OUT : out std_logic;  
            BYTE_LEN_OUT : out std_logic_vector (1 downto 0);  WB_LATCH_EN, 
            JAL_MUX_SEL, WB_MUX_SEL : in std_logic;  IR_IN : in 
            std_logic_vector (31 downto 0);  PC_OUT : out std_logic_vector (31 
            downto 0);  MEM_DATA_OUT_INT : in std_logic_vector (31 downto 0);  
            MEM_ADDR_OUT, MEM_DATA_IN_PRIME : out std_logic_vector (31 downto 
            0));
   end component;
   
   signal IF_LATCH_EN, PC_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, 
      WR_EN, ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN
      , ALU_OPCODE_6_port, ALU_OPCODE_5_port, ALU_OPCODE_4_port, 
      ALU_OPCODE_3_port, ALU_OPCODE_2_port, ALU_OPCODE_1_port, 
      ALU_OPCODE_0_port, MEM_OUTREG_EN, ZERO_PADDING4, MEM_OUT_SEL, 
      BYTE_LEN_INT_1_port, BYTE_LEN_INT_0_port, DRAM_WE_INT, WB_LATCH_EN, 
      JAL_MUX_SEL, WB_MUX_SEL, IR_IN_31_port, IR_IN_30_port, IR_IN_29_port, 
      IR_IN_28_port, IR_IN_27_port, IR_IN_26_port, IR_IN_25_port, IR_IN_24_port
      , IR_IN_23_port, IR_IN_22_port, IR_IN_21_port, IR_IN_20_port, 
      IR_IN_19_port, IR_IN_18_port, IR_IN_17_port, IR_IN_16_port, IR_IN_15_port
      , IR_IN_14_port, IR_IN_13_port, IR_IN_12_port, IR_IN_11_port, 
      IR_IN_10_port, IR_IN_9_port, IR_IN_8_port, IR_IN_7_port, IR_IN_6_port, 
      IR_IN_5_port, IR_IN_4_port, IR_IN_3_port, IR_IN_2_port, IR_IN_1_port, 
      IR_IN_0_port, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, 
      n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, 
      n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, 
      n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, 
      n_2246, n_2247, n_2248 : std_logic;

begin
   
   DATAPATH : 
                           DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 
                           port map( CLK => Clock, RST => ResetN, IF_LATCH_EN 
                           => IF_LATCH_EN, PC_LATCH_EN => PC_LATCH_EN, 
                           DEC_OUTREG_EN => DEC_OUTREG_EN, IS_I_TYPE => 
                           IS_I_TYPE, RD1_EN => RD1_EN, RD2_EN => RD2_EN, WR_EN
                           => WR_EN, ZERO_PADDING2 => ZERO_PADDING2, MUXA_SEL 
                           => MUXA_SEL, MUXB_SEL => MUXB_SEL, EXE_OUTREG_EN => 
                           EXE_OUTREG_EN, EQ_COND => EQ_COND, JUMP_EN => 
                           JUMP_EN, ALU_OPCODE(0) => ALU_OPCODE_6_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_5_port, ALU_OPCODE(2) =>
                           ALU_OPCODE_4_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_2_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_1_port, ALU_OPCODE(6) => 
                           ALU_OPCODE_0_port, MEM_OUTREG_EN => MEM_OUTREG_EN, 
                           ZERO_PADDING4 => ZERO_PADDING4, MEM_OUT_SEL => 
                           MEM_OUT_SEL, BYTE_LEN_IN(1) => BYTE_LEN_INT_1_port, 
                           BYTE_LEN_IN(0) => BYTE_LEN_INT_0_port, DRAM_WE => 
                           DRAM_WE_INT, DRAM_WE_OUT => DataMem_WrEn, 
                           BYTE_LEN_OUT(1) => DataMem_BLen(1), BYTE_LEN_OUT(0) 
                           => DataMem_BLen(0), WB_LATCH_EN => WB_LATCH_EN, 
                           JAL_MUX_SEL => JAL_MUX_SEL, WB_MUX_SEL => WB_MUX_SEL
                           , IR_IN(31) => IR_IN_31_port, IR_IN(30) => 
                           IR_IN_30_port, IR_IN(29) => IR_IN_29_port, IR_IN(28)
                           => IR_IN_28_port, IR_IN(27) => IR_IN_27_port, 
                           IR_IN(26) => IR_IN_26_port, IR_IN(25) => 
                           IR_IN_25_port, IR_IN(24) => IR_IN_24_port, IR_IN(23)
                           => IR_IN_23_port, IR_IN(22) => IR_IN_22_port, 
                           IR_IN(21) => IR_IN_21_port, IR_IN(20) => 
                           IR_IN_20_port, IR_IN(19) => IR_IN_19_port, IR_IN(18)
                           => IR_IN_18_port, IR_IN(17) => IR_IN_17_port, 
                           IR_IN(16) => IR_IN_16_port, IR_IN(15) => 
                           IR_IN_15_port, IR_IN(14) => IR_IN_14_port, IR_IN(13)
                           => IR_IN_13_port, IR_IN(12) => IR_IN_12_port, 
                           IR_IN(11) => IR_IN_11_port, IR_IN(10) => 
                           IR_IN_10_port, IR_IN(9) => IR_IN_9_port, IR_IN(8) =>
                           IR_IN_8_port, IR_IN(7) => IR_IN_7_port, IR_IN(6) => 
                           IR_IN_6_port, IR_IN(5) => IR_IN_5_port, IR_IN(4) => 
                           IR_IN_4_port, IR_IN(3) => IR_IN_3_port, IR_IN(2) => 
                           IR_IN_2_port, IR_IN(1) => IR_IN_1_port, IR_IN(0) => 
                           IR_IN_0_port, PC_OUT(31) => ProgCount_Out(31), 
                           PC_OUT(30) => ProgCount_Out(30), PC_OUT(29) => 
                           ProgCount_Out(29), PC_OUT(28) => ProgCount_Out(28), 
                           PC_OUT(27) => ProgCount_Out(27), PC_OUT(26) => 
                           ProgCount_Out(26), PC_OUT(25) => ProgCount_Out(25), 
                           PC_OUT(24) => ProgCount_Out(24), PC_OUT(23) => 
                           ProgCount_Out(23), PC_OUT(22) => ProgCount_Out(22), 
                           PC_OUT(21) => ProgCount_Out(21), PC_OUT(20) => 
                           ProgCount_Out(20), PC_OUT(19) => ProgCount_Out(19), 
                           PC_OUT(18) => ProgCount_Out(18), PC_OUT(17) => 
                           ProgCount_Out(17), PC_OUT(16) => ProgCount_Out(16), 
                           PC_OUT(15) => ProgCount_Out(15), PC_OUT(14) => 
                           ProgCount_Out(14), PC_OUT(13) => ProgCount_Out(13), 
                           PC_OUT(12) => ProgCount_Out(12), PC_OUT(11) => 
                           ProgCount_Out(11), PC_OUT(10) => ProgCount_Out(10), 
                           PC_OUT(9) => ProgCount_Out(9), PC_OUT(8) => 
                           ProgCount_Out(8), PC_OUT(7) => ProgCount_Out(7), 
                           PC_OUT(6) => ProgCount_Out(6), PC_OUT(5) => 
                           ProgCount_Out(5), PC_OUT(4) => ProgCount_Out(4), 
                           PC_OUT(3) => ProgCount_Out(3), PC_OUT(2) => 
                           ProgCount_Out(2), PC_OUT(1) => ProgCount_Out(1), 
                           PC_OUT(0) => ProgCount_Out(0), MEM_DATA_OUT_INT(31) 
                           => DataMem_Read(31), MEM_DATA_OUT_INT(30) => 
                           DataMem_Read(30), MEM_DATA_OUT_INT(29) => 
                           DataMem_Read(29), MEM_DATA_OUT_INT(28) => 
                           DataMem_Read(28), MEM_DATA_OUT_INT(27) => 
                           DataMem_Read(27), MEM_DATA_OUT_INT(26) => 
                           DataMem_Read(26), MEM_DATA_OUT_INT(25) => 
                           DataMem_Read(25), MEM_DATA_OUT_INT(24) => 
                           DataMem_Read(24), MEM_DATA_OUT_INT(23) => 
                           DataMem_Read(23), MEM_DATA_OUT_INT(22) => 
                           DataMem_Read(22), MEM_DATA_OUT_INT(21) => 
                           DataMem_Read(21), MEM_DATA_OUT_INT(20) => 
                           DataMem_Read(20), MEM_DATA_OUT_INT(19) => 
                           DataMem_Read(19), MEM_DATA_OUT_INT(18) => 
                           DataMem_Read(18), MEM_DATA_OUT_INT(17) => 
                           DataMem_Read(17), MEM_DATA_OUT_INT(16) => 
                           DataMem_Read(16), MEM_DATA_OUT_INT(15) => 
                           DataMem_Read(15), MEM_DATA_OUT_INT(14) => 
                           DataMem_Read(14), MEM_DATA_OUT_INT(13) => 
                           DataMem_Read(13), MEM_DATA_OUT_INT(12) => 
                           DataMem_Read(12), MEM_DATA_OUT_INT(11) => 
                           DataMem_Read(11), MEM_DATA_OUT_INT(10) => 
                           DataMem_Read(10), MEM_DATA_OUT_INT(9) => 
                           DataMem_Read(9), MEM_DATA_OUT_INT(8) => 
                           DataMem_Read(8), MEM_DATA_OUT_INT(7) => 
                           DataMem_Read(7), MEM_DATA_OUT_INT(6) => 
                           DataMem_Read(6), MEM_DATA_OUT_INT(5) => 
                           DataMem_Read(5), MEM_DATA_OUT_INT(4) => 
                           DataMem_Read(4), MEM_DATA_OUT_INT(3) => 
                           DataMem_Read(3), MEM_DATA_OUT_INT(2) => 
                           DataMem_Read(2), MEM_DATA_OUT_INT(1) => 
                           DataMem_Read(1), MEM_DATA_OUT_INT(0) => 
                           DataMem_Read(0), MEM_ADDR_OUT(31) => 
                           DataMem_Addr(31), MEM_ADDR_OUT(30) => 
                           DataMem_Addr(30), MEM_ADDR_OUT(29) => 
                           DataMem_Addr(29), MEM_ADDR_OUT(28) => 
                           DataMem_Addr(28), MEM_ADDR_OUT(27) => 
                           DataMem_Addr(27), MEM_ADDR_OUT(26) => 
                           DataMem_Addr(26), MEM_ADDR_OUT(25) => 
                           DataMem_Addr(25), MEM_ADDR_OUT(24) => 
                           DataMem_Addr(24), MEM_ADDR_OUT(23) => 
                           DataMem_Addr(23), MEM_ADDR_OUT(22) => 
                           DataMem_Addr(22), MEM_ADDR_OUT(21) => 
                           DataMem_Addr(21), MEM_ADDR_OUT(20) => 
                           DataMem_Addr(20), MEM_ADDR_OUT(19) => 
                           DataMem_Addr(19), MEM_ADDR_OUT(18) => 
                           DataMem_Addr(18), MEM_ADDR_OUT(17) => 
                           DataMem_Addr(17), MEM_ADDR_OUT(16) => 
                           DataMem_Addr(16), MEM_ADDR_OUT(15) => 
                           DataMem_Addr(15), MEM_ADDR_OUT(14) => 
                           DataMem_Addr(14), MEM_ADDR_OUT(13) => 
                           DataMem_Addr(13), MEM_ADDR_OUT(12) => 
                           DataMem_Addr(12), MEM_ADDR_OUT(11) => 
                           DataMem_Addr(11), MEM_ADDR_OUT(10) => 
                           DataMem_Addr(10), MEM_ADDR_OUT(9) => DataMem_Addr(9)
                           , MEM_ADDR_OUT(8) => DataMem_Addr(8), 
                           MEM_ADDR_OUT(7) => DataMem_Addr(7), MEM_ADDR_OUT(6) 
                           => DataMem_Addr(6), MEM_ADDR_OUT(5) => 
                           DataMem_Addr(5), MEM_ADDR_OUT(4) => DataMem_Addr(4),
                           MEM_ADDR_OUT(3) => DataMem_Addr(3), MEM_ADDR_OUT(2) 
                           => DataMem_Addr(2), MEM_ADDR_OUT(1) => 
                           DataMem_Addr(1), MEM_ADDR_OUT(0) => DataMem_Addr(0),
                           MEM_DATA_IN_PRIME(31) => DataMem_Write(31), 
                           MEM_DATA_IN_PRIME(30) => DataMem_Write(30), 
                           MEM_DATA_IN_PRIME(29) => DataMem_Write(29), 
                           MEM_DATA_IN_PRIME(28) => DataMem_Write(28), 
                           MEM_DATA_IN_PRIME(27) => DataMem_Write(27), 
                           MEM_DATA_IN_PRIME(26) => DataMem_Write(26), 
                           MEM_DATA_IN_PRIME(25) => DataMem_Write(25), 
                           MEM_DATA_IN_PRIME(24) => DataMem_Write(24), 
                           MEM_DATA_IN_PRIME(23) => DataMem_Write(23), 
                           MEM_DATA_IN_PRIME(22) => DataMem_Write(22), 
                           MEM_DATA_IN_PRIME(21) => DataMem_Write(21), 
                           MEM_DATA_IN_PRIME(20) => DataMem_Write(20), 
                           MEM_DATA_IN_PRIME(19) => DataMem_Write(19), 
                           MEM_DATA_IN_PRIME(18) => DataMem_Write(18), 
                           MEM_DATA_IN_PRIME(17) => DataMem_Write(17), 
                           MEM_DATA_IN_PRIME(16) => DataMem_Write(16), 
                           MEM_DATA_IN_PRIME(15) => DataMem_Write(15), 
                           MEM_DATA_IN_PRIME(14) => DataMem_Write(14), 
                           MEM_DATA_IN_PRIME(13) => DataMem_Write(13), 
                           MEM_DATA_IN_PRIME(12) => DataMem_Write(12), 
                           MEM_DATA_IN_PRIME(11) => DataMem_Write(11), 
                           MEM_DATA_IN_PRIME(10) => DataMem_Write(10), 
                           MEM_DATA_IN_PRIME(9) => DataMem_Write(9), 
                           MEM_DATA_IN_PRIME(8) => DataMem_Write(8), 
                           MEM_DATA_IN_PRIME(7) => DataMem_Write(7), 
                           MEM_DATA_IN_PRIME(6) => DataMem_Write(6), 
                           MEM_DATA_IN_PRIME(5) => DataMem_Write(5), 
                           MEM_DATA_IN_PRIME(4) => DataMem_Write(4), 
                           MEM_DATA_IN_PRIME(3) => DataMem_Write(3), 
                           MEM_DATA_IN_PRIME(2) => DataMem_Write(2), 
                           MEM_DATA_IN_PRIME(1) => DataMem_Write(1), 
                           MEM_DATA_IN_PRIME(0) => DataMem_Write(0));
   CONTROL : CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE22 
                           port map( Clk => Clock, Rst => ResetN, IR_IN(31) => 
                           Instr_In(31), IR_IN(30) => Instr_In(30), IR_IN(29) 
                           => Instr_In(29), IR_IN(28) => Instr_In(28), 
                           IR_IN(27) => Instr_In(27), IR_IN(26) => Instr_In(26)
                           , IR_IN(25) => Instr_In(25), IR_IN(24) => 
                           Instr_In(24), IR_IN(23) => Instr_In(23), IR_IN(22) 
                           => Instr_In(22), IR_IN(21) => Instr_In(21), 
                           IR_IN(20) => Instr_In(20), IR_IN(19) => Instr_In(19)
                           , IR_IN(18) => Instr_In(18), IR_IN(17) => 
                           Instr_In(17), IR_IN(16) => Instr_In(16), IR_IN(15) 
                           => Instr_In(15), IR_IN(14) => Instr_In(14), 
                           IR_IN(13) => Instr_In(13), IR_IN(12) => Instr_In(12)
                           , IR_IN(11) => Instr_In(11), IR_IN(10) => 
                           Instr_In(10), IR_IN(9) => Instr_In(9), IR_IN(8) => 
                           Instr_In(8), IR_IN(7) => Instr_In(7), IR_IN(6) => 
                           Instr_In(6), IR_IN(5) => Instr_In(5), IR_IN(4) => 
                           Instr_In(4), IR_IN(3) => Instr_In(3), IR_IN(2) => 
                           Instr_In(2), IR_IN(1) => Instr_In(1), IR_IN(0) => 
                           Instr_In(0), IF_LATCH_EN => IF_LATCH_EN, 
                           DEC_OUTREG_EN => DEC_OUTREG_EN, IS_I_TYPE => 
                           IS_I_TYPE, RD1_EN => RD1_EN, RD2_EN => RD2_EN, 
                           ZERO_PADDING2 => ZERO_PADDING2, MUXA_SEL => MUXA_SEL
                           , MUXB_SEL => MUXB_SEL, EXE_OUTREG_EN => 
                           EXE_OUTREG_EN, EQ_COND => EQ_COND, JUMP_EN => 
                           JUMP_EN, ALU_OPCODE(0) => ALU_OPCODE_6_port, 
                           ALU_OPCODE(1) => ALU_OPCODE_5_port, ALU_OPCODE(2) =>
                           ALU_OPCODE_4_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_3_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_2_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_1_port, ALU_OPCODE(6) => 
                           ALU_OPCODE_0_port, FPU_OPCODE(0) => n_2212, 
                           FPU_OPCODE(1) => n_2213, FPU_OPCODE(2) => n_2214, 
                           FPU_OPCODE(3) => n_2215, FPU_OPCODE(4) => n_2216, 
                           PC_LATCH_EN => PC_LATCH_EN, MEM_OUTREG_EN => 
                           MEM_OUTREG_EN, ZERO_PADDING4 => ZERO_PADDING4, 
                           MEM_OUT_SEL => MEM_OUT_SEL, DRAM_WE => DRAM_WE_INT, 
                           BYTE_LEN(1) => BYTE_LEN_INT_1_port, BYTE_LEN(0) => 
                           BYTE_LEN_INT_0_port, WB_MUX_SEL => WB_MUX_SEL, 
                           JAL_MUX_SEL => JAL_MUX_SEL, WR_EN => WR_EN, 
                           WB_LATCH_EN => WB_LATCH_EN);
   IR_IN_reg_31_inst : DFFR_X1 port map( D => Instr_In(31), CK => Clock, RN => 
                           ResetN, Q => IR_IN_31_port, QN => n_2217);
   IR_IN_reg_30_inst : DFFR_X1 port map( D => Instr_In(30), CK => Clock, RN => 
                           ResetN, Q => IR_IN_30_port, QN => n_2218);
   IR_IN_reg_29_inst : DFFR_X1 port map( D => Instr_In(29), CK => Clock, RN => 
                           ResetN, Q => IR_IN_29_port, QN => n_2219);
   IR_IN_reg_28_inst : DFFR_X1 port map( D => Instr_In(28), CK => Clock, RN => 
                           ResetN, Q => IR_IN_28_port, QN => n_2220);
   IR_IN_reg_27_inst : DFFR_X1 port map( D => Instr_In(27), CK => Clock, RN => 
                           ResetN, Q => IR_IN_27_port, QN => n_2221);
   IR_IN_reg_26_inst : DFFR_X1 port map( D => Instr_In(26), CK => Clock, RN => 
                           ResetN, Q => IR_IN_26_port, QN => n_2222);
   IR_IN_reg_25_inst : DFFR_X1 port map( D => Instr_In(25), CK => Clock, RN => 
                           ResetN, Q => IR_IN_25_port, QN => n_2223);
   IR_IN_reg_24_inst : DFFR_X1 port map( D => Instr_In(24), CK => Clock, RN => 
                           ResetN, Q => IR_IN_24_port, QN => n_2224);
   IR_IN_reg_23_inst : DFFR_X1 port map( D => Instr_In(23), CK => Clock, RN => 
                           ResetN, Q => IR_IN_23_port, QN => n_2225);
   IR_IN_reg_22_inst : DFFR_X1 port map( D => Instr_In(22), CK => Clock, RN => 
                           ResetN, Q => IR_IN_22_port, QN => n_2226);
   IR_IN_reg_21_inst : DFFR_X1 port map( D => Instr_In(21), CK => Clock, RN => 
                           ResetN, Q => IR_IN_21_port, QN => n_2227);
   IR_IN_reg_20_inst : DFFR_X1 port map( D => Instr_In(20), CK => Clock, RN => 
                           ResetN, Q => IR_IN_20_port, QN => n_2228);
   IR_IN_reg_19_inst : DFFR_X1 port map( D => Instr_In(19), CK => Clock, RN => 
                           ResetN, Q => IR_IN_19_port, QN => n_2229);
   IR_IN_reg_18_inst : DFFR_X1 port map( D => Instr_In(18), CK => Clock, RN => 
                           ResetN, Q => IR_IN_18_port, QN => n_2230);
   IR_IN_reg_17_inst : DFFR_X1 port map( D => Instr_In(17), CK => Clock, RN => 
                           ResetN, Q => IR_IN_17_port, QN => n_2231);
   IR_IN_reg_16_inst : DFFR_X1 port map( D => Instr_In(16), CK => Clock, RN => 
                           ResetN, Q => IR_IN_16_port, QN => n_2232);
   IR_IN_reg_15_inst : DFFR_X1 port map( D => Instr_In(15), CK => Clock, RN => 
                           ResetN, Q => IR_IN_15_port, QN => n_2233);
   IR_IN_reg_14_inst : DFFR_X1 port map( D => Instr_In(14), CK => Clock, RN => 
                           ResetN, Q => IR_IN_14_port, QN => n_2234);
   IR_IN_reg_13_inst : DFFR_X1 port map( D => Instr_In(13), CK => Clock, RN => 
                           ResetN, Q => IR_IN_13_port, QN => n_2235);
   IR_IN_reg_12_inst : DFFR_X1 port map( D => Instr_In(12), CK => Clock, RN => 
                           ResetN, Q => IR_IN_12_port, QN => n_2236);
   IR_IN_reg_11_inst : DFFR_X1 port map( D => Instr_In(11), CK => Clock, RN => 
                           ResetN, Q => IR_IN_11_port, QN => n_2237);
   IR_IN_reg_10_inst : DFFR_X1 port map( D => Instr_In(10), CK => Clock, RN => 
                           ResetN, Q => IR_IN_10_port, QN => n_2238);
   IR_IN_reg_9_inst : DFFR_X1 port map( D => Instr_In(9), CK => Clock, RN => 
                           ResetN, Q => IR_IN_9_port, QN => n_2239);
   IR_IN_reg_8_inst : DFFR_X1 port map( D => Instr_In(8), CK => Clock, RN => 
                           ResetN, Q => IR_IN_8_port, QN => n_2240);
   IR_IN_reg_7_inst : DFFR_X1 port map( D => Instr_In(7), CK => Clock, RN => 
                           ResetN, Q => IR_IN_7_port, QN => n_2241);
   IR_IN_reg_6_inst : DFFR_X1 port map( D => Instr_In(6), CK => Clock, RN => 
                           ResetN, Q => IR_IN_6_port, QN => n_2242);
   IR_IN_reg_5_inst : DFFR_X1 port map( D => Instr_In(5), CK => Clock, RN => 
                           ResetN, Q => IR_IN_5_port, QN => n_2243);
   IR_IN_reg_4_inst : DFFR_X1 port map( D => Instr_In(4), CK => Clock, RN => 
                           ResetN, Q => IR_IN_4_port, QN => n_2244);
   IR_IN_reg_3_inst : DFFR_X1 port map( D => Instr_In(3), CK => Clock, RN => 
                           ResetN, Q => IR_IN_3_port, QN => n_2245);
   IR_IN_reg_2_inst : DFFR_X1 port map( D => Instr_In(2), CK => Clock, RN => 
                           ResetN, Q => IR_IN_2_port, QN => n_2246);
   IR_IN_reg_1_inst : DFFR_X1 port map( D => Instr_In(1), CK => Clock, RN => 
                           ResetN, Q => IR_IN_1_port, QN => n_2247);
   IR_IN_reg_0_inst : DFFR_X1 port map( D => Instr_In(0), CK => Clock, RN => 
                           ResetN, Q => IR_IN_0_port, QN => n_2248);

end SYN_PRO;
