
module gen_reg_N32_0 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, net76207, net76206,
         net76215, net76214, net82947, n70, net82630, net74891, n69, n97;

  DFFR_X2 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[30]), 
        .QN(n2) );
  OAI21_X1 U2 ( .B1(n38), .B2(n97), .A(n65), .ZN(n9) );
  NAND2_X1 U3 ( .A1(net76215), .A2(data_in[26]), .ZN(n65) );
  OAI21_X1 U4 ( .B1(n37), .B2(net76207), .A(n66), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(net76214), .ZN(n66) );
  OAI21_X1 U6 ( .B1(n36), .B2(n97), .A(n67), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(net76214), .ZN(n67) );
  OAI21_X1 U8 ( .B1(n3), .B2(n97), .A(n68), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(net76214), .ZN(n68) );
  OAI21_X1 U14 ( .B1(n64), .B2(net76206), .A(n71), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(net76214), .ZN(n71) );
  OAI21_X1 U16 ( .B1(n63), .B2(net74891), .A(n72), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(net76215), .ZN(n72) );
  OAI21_X1 U18 ( .B1(n62), .B2(net76207), .A(n73), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(net76215), .ZN(n73) );
  OAI21_X1 U20 ( .B1(n61), .B2(n97), .A(n74), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(net76215), .ZN(n74) );
  OAI21_X1 U22 ( .B1(n60), .B2(net74891), .A(n75), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(net74891), .ZN(n75) );
  OAI21_X1 U24 ( .B1(n59), .B2(net76215), .A(n76), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n97), .ZN(n76) );
  OAI21_X1 U26 ( .B1(n58), .B2(net76214), .A(n77), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(ld), .ZN(n77) );
  OAI21_X1 U28 ( .B1(n57), .B2(n97), .A(n78), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n97), .ZN(n78) );
  OAI21_X1 U30 ( .B1(n56), .B2(net76207), .A(n79), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(net74891), .ZN(n79) );
  OAI21_X1 U32 ( .B1(n55), .B2(net74891), .A(n80), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(net74891), .ZN(n80) );
  OAI21_X1 U34 ( .B1(n54), .B2(net76207), .A(n81), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(n97), .ZN(n81) );
  OAI21_X1 U36 ( .B1(n53), .B2(n97), .A(n82), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(net74891), .ZN(n82) );
  OAI21_X1 U38 ( .B1(n52), .B2(net76207), .A(n83), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(ld), .ZN(n83) );
  OAI21_X1 U40 ( .B1(n51), .B2(net76207), .A(n84), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(net74891), .ZN(n84) );
  OAI21_X1 U42 ( .B1(n50), .B2(net76206), .A(n85), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(net74891), .ZN(n85) );
  OAI21_X1 U44 ( .B1(n49), .B2(net76207), .A(n86), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(net74891), .ZN(n86) );
  OAI21_X1 U46 ( .B1(n48), .B2(net76207), .A(n87), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n97), .ZN(n87) );
  OAI21_X1 U48 ( .B1(n47), .B2(net76207), .A(n88), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n97), .ZN(n88) );
  OAI21_X1 U50 ( .B1(n46), .B2(net76207), .A(n89), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(net74891), .ZN(n89) );
  OAI21_X1 U52 ( .B1(n45), .B2(net76206), .A(n90), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(net74891), .ZN(n90) );
  OAI21_X1 U54 ( .B1(n44), .B2(net76206), .A(n91), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n97), .ZN(n91) );
  OAI21_X1 U56 ( .B1(n43), .B2(net74891), .A(n92), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(net74891), .ZN(n92) );
  OAI21_X1 U58 ( .B1(n42), .B2(net76206), .A(n93), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(n97), .ZN(n93) );
  OAI21_X1 U60 ( .B1(n41), .B2(n97), .A(n94), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(ld), .ZN(n94) );
  OAI21_X1 U62 ( .B1(n40), .B2(net74891), .A(n95), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n97), .ZN(n95) );
  OAI21_X1 U64 ( .B1(n39), .B2(n97), .A(n96), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(net74891), .ZN(n96) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(net76214), .ZN(n70) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(net76215), .ZN(n69) );
  NAND2_X1 U10 ( .A1(n69), .A2(net82630), .ZN(n5) );
  OR2_X1 U12 ( .A1(n2), .A2(net76206), .ZN(net82630) );
  CLKBUF_X1 U66 ( .A(net74891), .Z(net76206) );
  CLKBUF_X1 U67 ( .A(ld), .Z(net74891) );
  CLKBUF_X1 U68 ( .A(net74891), .Z(net76207) );
  CLKBUF_X1 U69 ( .A(n97), .Z(net76215) );
  CLKBUF_X1 U70 ( .A(ld), .Z(n97) );
  CLKBUF_X1 U71 ( .A(n97), .Z(net76214) );
  NAND2_X1 U72 ( .A1(n70), .A2(net82947), .ZN(n4) );
  OR2_X1 U73 ( .A1(n1), .A2(net76206), .ZN(net82947) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[31]), 
        .QN(n1) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(rst), .Q(data_out[29]), 
        .QN(n3) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(rst), .Q(data_out[28]), 
        .QN(n36) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(rst), .Q(data_out[27]), 
        .QN(n37) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(rst), .Q(data_out[26]), 
        .QN(n38) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(rst), .Q(data_out[25]), 
        .QN(n39) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(rst), .Q(data_out[24]), 
        .QN(n40) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(rst), .Q(data_out[23]), 
        .QN(n41) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(rst), .Q(data_out[22]), 
        .QN(n42) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(rst), .Q(data_out[21]), 
        .QN(n43) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(rst), .Q(data_out[20]), 
        .QN(n44) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(rst), .Q(data_out[19]), 
        .QN(n45) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(rst), .Q(data_out[18]), 
        .QN(n46) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n47) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n48) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n49) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n50) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n51) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(rst), .Q(data_out[12]), 
        .QN(n52) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(rst), .Q(data_out[11]), 
        .QN(n53) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(rst), .Q(data_out[10]), 
        .QN(n54) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(rst), .Q(data_out[9]), 
        .QN(n55) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(rst), .Q(data_out[8]), 
        .QN(n56) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(rst), .Q(data_out[7]), 
        .QN(n57) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(rst), .Q(data_out[6]), 
        .QN(n58) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(rst), .Q(data_out[5]), 
        .QN(n59) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n60) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n61) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n62) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n63) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n64) );
endmodule


module gen_reg_N32_11 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n97, n98, n112, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181;

  OAI21_X1 U2 ( .B1(n176), .B2(n112), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n97), .A2(data_in[26]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n177), .B2(ld), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(n112), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n178), .B2(n112), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(n97), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n179), .B2(ld), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(n97), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n180), .B2(n112), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(n112), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n181), .B2(n112), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(n97), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n98), .A(n143), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n112), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n98), .A(n142), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n112), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n98), .A(n141), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n97), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n153), .B2(n98), .A(n140), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(n112), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n154), .B2(n98), .A(n139), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(n97), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n155), .B2(n112), .A(n138), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n97), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n156), .B2(n98), .A(n137), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(n112), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n157), .B2(n98), .A(n136), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n97), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n158), .B2(n98), .A(n135), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(n97), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n159), .B2(n98), .A(n134), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(n97), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n160), .B2(n98), .A(n133), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(n97), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n161), .B2(n98), .A(n132), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(n97), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n162), .B2(n112), .A(n131), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(n97), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n163), .B2(n98), .A(n130), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(n97), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n164), .B2(n112), .A(n129), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(n97), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n165), .B2(n112), .A(n128), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(n98), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n166), .B2(n97), .A(n127), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n97), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n167), .B2(n112), .A(n126), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n98), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n168), .B2(n112), .A(n125), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(n97), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n169), .B2(n112), .A(n124), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(n98), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n170), .B2(n97), .A(n123), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n97), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n171), .B2(n97), .A(n122), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(n98), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n172), .B2(n112), .A(n121), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(n97), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n173), .B2(n98), .A(n120), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(n98), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n174), .B2(n112), .A(n119), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n97), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n175), .B2(n112), .A(n118), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(n97), .ZN(n118) );
  CLKBUF_X1 U69 ( .A(ld), .Z(n97) );
  CLKBUF_X1 U75 ( .A(ld), .Z(n98) );
  CLKBUF_X1 U84 ( .A(ld), .Z(n112) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(rst), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(rst), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(rst), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(rst), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(rst), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(rst), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(rst), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(rst), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(rst), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(rst), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(rst), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(rst), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(rst), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(rst), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(rst), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(rst), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(rst), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(rst), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(rst), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(rst), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N32_10 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n101, n102, n110, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n176), .B2(n101), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n102), .A2(data_in[26]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n177), .B2(n102), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(n101), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n178), .B2(ld), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(n101), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n179), .B2(n101), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(n101), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n180), .B2(n110), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(n102), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n181), .B2(n110), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(n101), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n102), .A(n143), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n101), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n102), .A(n142), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n102), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n102), .A(n141), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n102), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n153), .B2(n110), .A(n140), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(n102), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n154), .B2(n110), .A(n139), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(n110), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n155), .B2(n102), .A(n138), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n110), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n156), .B2(n110), .A(n137), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(n110), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n157), .B2(n102), .A(n136), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n110), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n158), .B2(n102), .A(n135), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(n110), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n159), .B2(n102), .A(n134), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(n102), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n160), .B2(ld), .A(n133), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(n110), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n161), .B2(n101), .A(n132), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(n101), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n162), .B2(ld), .A(n131), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(n110), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n163), .B2(ld), .A(n130), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(n101), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n164), .B2(n101), .A(n129), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(n110), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n165), .B2(ld), .A(n128), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(n101), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n166), .B2(n110), .A(n127), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n110), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n167), .B2(n101), .A(n126), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n102), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n168), .B2(n102), .A(n125), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(n101), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n169), .B2(n102), .A(n124), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(n102), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n170), .B2(ld), .A(n123), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n101), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n171), .B2(n101), .A(n122), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(n102), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n172), .B2(n101), .A(n121), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(ld), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n173), .B2(n101), .A(n120), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(n101), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n174), .B2(n101), .A(n119), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n102), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n175), .B2(n101), .A(n118), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(n102), .ZN(n118) );
  CLKBUF_X1 U67 ( .A(rst), .Z(n116) );
  CLKBUF_X1 U68 ( .A(rst), .Z(n117) );
  CLKBUF_X1 U71 ( .A(ld), .Z(n102) );
  CLKBUF_X1 U76 ( .A(ld), .Z(n101) );
  CLKBUF_X1 U82 ( .A(ld), .Z(n110) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(n117), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(n117), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(n117), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(n117), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(n117), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(n117), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(n117), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(n117), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(n117), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(n117), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(n116), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(n116), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(n116), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(n116), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(n116), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(n116), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(n116), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(n116), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(n116), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(n116), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(n116), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(n116), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(n117), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(n116), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(n117), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(n116), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(n117), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(n116), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(n117), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(n116), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(n117), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N32_9 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n99, n100, n110, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n176), .B2(n110), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n110), .A2(data_in[26]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n177), .B2(n99), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(n110), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n178), .B2(n100), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(ld), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n179), .B2(n99), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(n100), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n180), .B2(n110), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(n99), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n181), .B2(n99), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(n100), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n100), .A(n143), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n110), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n110), .A(n142), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n100), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n99), .A(n141), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n99), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n153), .B2(n110), .A(n140), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(n110), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n154), .B2(n110), .A(n139), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(n100), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n155), .B2(n110), .A(n138), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n99), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n156), .B2(n110), .A(n137), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(n100), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n157), .B2(n110), .A(n136), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n99), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n158), .B2(n100), .A(n135), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(n100), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n159), .B2(n100), .A(n134), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(n99), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n160), .B2(n110), .A(n133), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(n100), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n161), .B2(n110), .A(n132), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(n99), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n162), .B2(n99), .A(n131), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(n100), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n163), .B2(n100), .A(n130), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(n99), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n164), .B2(ld), .A(n129), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(n99), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n165), .B2(n110), .A(n128), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(n99), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n166), .B2(n100), .A(n127), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n100), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n167), .B2(n99), .A(n126), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n100), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n168), .B2(n100), .A(n125), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(n110), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n169), .B2(n110), .A(n124), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(n99), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n170), .B2(n99), .A(n123), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n110), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n171), .B2(n110), .A(n122), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(n99), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n172), .B2(n110), .A(n121), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(n110), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n173), .B2(n100), .A(n120), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(n110), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n174), .B2(n110), .A(n119), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n100), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n175), .B2(n100), .A(n118), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(n99), .ZN(n118) );
  CLKBUF_X1 U67 ( .A(rst), .Z(n116) );
  CLKBUF_X1 U68 ( .A(rst), .Z(n117) );
  CLKBUF_X1 U70 ( .A(n110), .Z(n99) );
  CLKBUF_X1 U74 ( .A(n110), .Z(n100) );
  CLKBUF_X1 U82 ( .A(ld), .Z(n110) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(n117), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(n117), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(n117), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(n117), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(n117), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(n117), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(n117), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(n117), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(n117), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(n117), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(n116), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(n116), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(n116), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(n116), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(n116), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(n116), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(n116), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(n116), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(n116), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(n116), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(n116), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(n116), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(n117), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(n116), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(n117), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(n116), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(n117), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(n116), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(n117), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N32_8 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n98, n99, n109, n115, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n176), .B2(n98), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n109), .A2(data_in[26]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n177), .B2(n98), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(n109), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n178), .B2(n98), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(n109), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n179), .B2(ld), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(n109), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n180), .B2(n98), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(n109), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n181), .B2(n99), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(n109), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n109), .A(n143), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n109), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n109), .A(n142), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n109), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n99), .A(n141), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n109), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n153), .B2(n109), .A(n140), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(n109), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n154), .B2(n98), .A(n139), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(n109), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n155), .B2(n109), .A(n138), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n99), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n156), .B2(n109), .A(n137), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(ld), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n157), .B2(n98), .A(n136), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n99), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n158), .B2(n109), .A(n135), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(n109), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n159), .B2(n109), .A(n134), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(n99), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n160), .B2(n99), .A(n133), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(ld), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n161), .B2(n98), .A(n132), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(n99), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n162), .B2(n98), .A(n131), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(n109), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n163), .B2(n109), .A(n130), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(n99), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n164), .B2(n109), .A(n129), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(n99), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n165), .B2(n99), .A(n128), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(n98), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n166), .B2(n98), .A(n127), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n98), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n167), .B2(n98), .A(n126), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n98), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n168), .B2(n99), .A(n125), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(n99), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n169), .B2(n98), .A(n124), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(n98), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n170), .B2(n109), .A(n123), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n99), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n171), .B2(n99), .A(n122), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(n98), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n172), .B2(n99), .A(n121), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(n99), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n173), .B2(n99), .A(n120), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(n98), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n174), .B2(ld), .A(n119), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n98), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n175), .B2(n98), .A(n118), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(n99), .ZN(n118) );
  CLKBUF_X1 U66 ( .A(rst), .Z(n115) );
  CLKBUF_X1 U70 ( .A(n109), .Z(n99) );
  CLKBUF_X1 U75 ( .A(n109), .Z(n98) );
  CLKBUF_X1 U81 ( .A(ld), .Z(n109) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(n115), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(n115), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(n115), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(n115), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(n115), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(n115), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(n115), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(n115), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(n115), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(n115), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(rst), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(rst), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(rst), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(rst), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(rst), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(rst), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(n115), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(n115), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(n115), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(n115), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(n115), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(n115), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(n115), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(n115), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(n115), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(n115), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(n115), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module pc_add_N32_OP24_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U29 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U30 ( .A(A[4]), .B(n1), .Z(SUM[4]) );
  XOR2_X1 U31 ( .A(A[5]), .B(n2), .Z(SUM[5]) );
  XOR2_X1 U32 ( .A(A[6]), .B(n3), .Z(SUM[6]) );
  XOR2_X1 U33 ( .A(A[7]), .B(n4), .Z(SUM[7]) );
  XOR2_X1 U34 ( .A(A[8]), .B(n5), .Z(SUM[8]) );
  XOR2_X1 U35 ( .A(A[9]), .B(n6), .Z(SUM[9]) );
  XOR2_X1 U36 ( .A(A[10]), .B(n7), .Z(SUM[10]) );
  XOR2_X1 U37 ( .A(A[11]), .B(n8), .Z(SUM[11]) );
  XOR2_X1 U38 ( .A(A[12]), .B(n9), .Z(SUM[12]) );
  XOR2_X1 U39 ( .A(A[13]), .B(n10), .Z(SUM[13]) );
  XOR2_X1 U40 ( .A(A[14]), .B(n11), .Z(SUM[14]) );
  XOR2_X1 U41 ( .A(A[15]), .B(n12), .Z(SUM[15]) );
  XOR2_X1 U42 ( .A(A[16]), .B(n13), .Z(SUM[16]) );
  XOR2_X1 U43 ( .A(A[17]), .B(n14), .Z(SUM[17]) );
  XOR2_X1 U44 ( .A(A[18]), .B(n15), .Z(SUM[18]) );
  XOR2_X1 U45 ( .A(A[19]), .B(n16), .Z(SUM[19]) );
  XOR2_X1 U46 ( .A(A[20]), .B(n17), .Z(SUM[20]) );
  XOR2_X1 U47 ( .A(A[21]), .B(n18), .Z(SUM[21]) );
  XOR2_X1 U48 ( .A(A[22]), .B(n19), .Z(SUM[22]) );
  XOR2_X1 U49 ( .A(A[23]), .B(n20), .Z(SUM[23]) );
  XOR2_X1 U50 ( .A(A[24]), .B(n21), .Z(SUM[24]) );
  XOR2_X1 U51 ( .A(A[25]), .B(n22), .Z(SUM[25]) );
  XOR2_X1 U52 ( .A(A[26]), .B(n23), .Z(SUM[26]) );
  XOR2_X1 U53 ( .A(A[27]), .B(n24), .Z(SUM[27]) );
  XOR2_X1 U54 ( .A(A[28]), .B(n25), .Z(SUM[28]) );
  XOR2_X1 U55 ( .A(A[29]), .B(n26), .Z(SUM[29]) );
  XOR2_X1 U56 ( .A(A[30]), .B(n27), .Z(SUM[30]) );
  XNOR2_X1 U57 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U58 ( .A1(A[30]), .A2(n27), .ZN(n57) );
  INV_X1 U28 ( .A(A[2]), .ZN(SUM[2]) );
  AND2_X1 U1 ( .A1(A[29]), .A2(n26), .ZN(n27) );
  AND2_X1 U2 ( .A1(A[3]), .A2(A[2]), .ZN(n1) );
  AND2_X1 U3 ( .A1(A[4]), .A2(n1), .ZN(n2) );
  AND2_X1 U4 ( .A1(A[5]), .A2(n2), .ZN(n3) );
  AND2_X1 U5 ( .A1(A[6]), .A2(n3), .ZN(n4) );
  AND2_X1 U6 ( .A1(A[7]), .A2(n4), .ZN(n5) );
  AND2_X1 U7 ( .A1(A[8]), .A2(n5), .ZN(n6) );
  AND2_X1 U8 ( .A1(A[9]), .A2(n6), .ZN(n7) );
  AND2_X1 U9 ( .A1(A[10]), .A2(n7), .ZN(n8) );
  AND2_X1 U10 ( .A1(A[11]), .A2(n8), .ZN(n9) );
  AND2_X1 U11 ( .A1(A[12]), .A2(n9), .ZN(n10) );
  AND2_X1 U12 ( .A1(A[13]), .A2(n10), .ZN(n11) );
  AND2_X1 U13 ( .A1(A[14]), .A2(n11), .ZN(n12) );
  AND2_X1 U14 ( .A1(A[15]), .A2(n12), .ZN(n13) );
  AND2_X1 U15 ( .A1(A[16]), .A2(n13), .ZN(n14) );
  AND2_X1 U16 ( .A1(A[17]), .A2(n14), .ZN(n15) );
  AND2_X1 U17 ( .A1(A[18]), .A2(n15), .ZN(n16) );
  AND2_X1 U18 ( .A1(A[19]), .A2(n16), .ZN(n17) );
  AND2_X1 U19 ( .A1(A[20]), .A2(n17), .ZN(n18) );
  AND2_X1 U20 ( .A1(A[21]), .A2(n18), .ZN(n19) );
  AND2_X1 U21 ( .A1(A[22]), .A2(n19), .ZN(n20) );
  AND2_X1 U22 ( .A1(A[23]), .A2(n20), .ZN(n21) );
  AND2_X1 U23 ( .A1(A[24]), .A2(n21), .ZN(n22) );
  AND2_X1 U24 ( .A1(A[25]), .A2(n22), .ZN(n23) );
  AND2_X1 U25 ( .A1(A[26]), .A2(n23), .ZN(n24) );
  AND2_X1 U26 ( .A1(A[27]), .A2(n24), .ZN(n25) );
  AND2_X1 U27 ( .A1(A[28]), .A2(n25), .ZN(n26) );
endmodule


module pc_add_N32_OP24 ( data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;


  pc_add_N32_OP24_DW01_add_0 add_21 ( .A(data_in), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(data_out) );
endmodule


module IF_STAGE_N_BITS_DATA32_N_BYTES_INST4 ( CLK, RST, IF_LATCH_EN, PC_IN, 
        IR_IN, PC_OUT, IR_OUT, ADD_OUT, NPC_OUT );
  input [31:0] PC_IN;
  input [31:0] IR_IN;
  output [31:0] PC_OUT;
  output [31:0] IR_OUT;
  output [31:0] ADD_OUT;
  output [31:0] NPC_OUT;
  input CLK, RST, IF_LATCH_EN;

  wire   [31:0] NPC_INTA;
  wire   [31:0] NPC_INTB;

  gen_reg_N32_0 PC ( .clk(CLK), .rst(RST), .ld(IF_LATCH_EN), .data_in(PC_IN), 
        .data_out(PC_OUT) );
  gen_reg_N32_11 IR ( .clk(CLK), .rst(RST), .ld(IF_LATCH_EN), .data_in(IR_IN), 
        .data_out(IR_OUT) );
  gen_reg_N32_10 NPC0 ( .clk(CLK), .rst(RST), .ld(IF_LATCH_EN), .data_in(
        ADD_OUT), .data_out(NPC_INTA) );
  gen_reg_N32_9 NPCA ( .clk(CLK), .rst(RST), .ld(IF_LATCH_EN), .data_in(
        NPC_INTA), .data_out(NPC_INTB) );
  gen_reg_N32_8 NPCB ( .clk(CLK), .rst(RST), .ld(IF_LATCH_EN), .data_in(
        NPC_INTB), .data_out(NPC_OUT) );
  pc_add_N32_OP24 PC_ADDER ( .data_in(PC_OUT), .data_out(ADD_OUT) );
endmodule


module gen_reg_N32_7 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n97, n98, n109, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n176), .B2(n97), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n109), .A2(data_in[26]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n177), .B2(n98), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(n109), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n178), .B2(n109), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(n97), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n179), .B2(n98), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(n109), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n180), .B2(n98), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(n98), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n181), .B2(n97), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(n109), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n98), .A(n143), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n97), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n97), .A(n142), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n109), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n98), .A(n141), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n109), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n153), .B2(n97), .A(n140), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(n109), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n154), .B2(n109), .A(n139), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(n97), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n155), .B2(n97), .A(n138), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n109), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n156), .B2(n109), .A(n137), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(n109), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n157), .B2(n109), .A(n136), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n98), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n158), .B2(n109), .A(n135), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(ld), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n159), .B2(n109), .A(n134), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(n109), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n160), .B2(n109), .A(n133), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(n109), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n161), .B2(n98), .A(n132), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(n109), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n162), .B2(n98), .A(n131), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(n109), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n163), .B2(n97), .A(n130), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(n98), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n164), .B2(n97), .A(n129), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(n97), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n165), .B2(n109), .A(n128), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(n98), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n166), .B2(n98), .A(n127), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n97), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n167), .B2(n109), .A(n126), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n98), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n168), .B2(ld), .A(n125), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(n97), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n169), .B2(ld), .A(n124), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(n98), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n170), .B2(n97), .A(n123), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n97), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n171), .B2(n98), .A(n122), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(n98), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n172), .B2(n98), .A(n121), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(n97), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n173), .B2(n97), .A(n120), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(n98), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n174), .B2(n98), .A(n119), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n97), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n175), .B2(n109), .A(n118), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(n97), .ZN(n118) );
  CLKBUF_X1 U67 ( .A(rst), .Z(n116) );
  CLKBUF_X1 U68 ( .A(rst), .Z(n117) );
  CLKBUF_X1 U69 ( .A(n109), .Z(n97) );
  CLKBUF_X1 U75 ( .A(n109), .Z(n98) );
  CLKBUF_X1 U81 ( .A(ld), .Z(n109) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(n117), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(n117), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(n117), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(n117), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(n117), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(n117), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(n117), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(n117), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(n117), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(n117), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(n116), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(n116), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(n116), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(n116), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(n116), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(n116), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(n116), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(n116), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(n116), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(n116), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(n116), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(n116), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(n117), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(n116), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(n117), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(n116), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(n117), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(n116), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(n117), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(n116), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(n117), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N32_6 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n99, n100, n109, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n176), .B2(ld), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n100), .A2(data_in[26]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n177), .B2(ld), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[27]), .A2(n99), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n178), .B2(n100), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[28]), .A2(n100), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n179), .B2(n99), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[29]), .A2(n99), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n180), .B2(n100), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[30]), .A2(n100), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n181), .B2(n99), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[31]), .A2(n100), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(ld), .A(n143), .ZN(n35) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n109), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n109), .A(n142), .ZN(n34) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n99), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n100), .A(n141), .ZN(n33) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n100), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n153), .B2(ld), .A(n140), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data_in[3]), .A2(n99), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n154), .B2(n100), .A(n139), .ZN(n31) );
  NAND2_X1 U23 ( .A1(data_in[4]), .A2(n100), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n155), .B2(n99), .A(n138), .ZN(n30) );
  NAND2_X1 U25 ( .A1(data_in[5]), .A2(n99), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n156), .B2(ld), .A(n137), .ZN(n29) );
  NAND2_X1 U27 ( .A1(data_in[6]), .A2(n100), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n157), .B2(ld), .A(n136), .ZN(n28) );
  NAND2_X1 U29 ( .A1(data_in[7]), .A2(n99), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n158), .B2(n109), .A(n135), .ZN(n27) );
  NAND2_X1 U31 ( .A1(data_in[8]), .A2(n100), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n159), .B2(n109), .A(n134), .ZN(n26) );
  NAND2_X1 U33 ( .A1(data_in[9]), .A2(n99), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n160), .B2(n109), .A(n133), .ZN(n25) );
  NAND2_X1 U35 ( .A1(data_in[10]), .A2(n100), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n161), .B2(n100), .A(n132), .ZN(n24) );
  NAND2_X1 U37 ( .A1(data_in[11]), .A2(n99), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n162), .B2(n100), .A(n131), .ZN(n23) );
  NAND2_X1 U39 ( .A1(data_in[12]), .A2(n100), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n163), .B2(ld), .A(n130), .ZN(n22) );
  NAND2_X1 U41 ( .A1(data_in[13]), .A2(n99), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n164), .B2(n99), .A(n129), .ZN(n21) );
  NAND2_X1 U43 ( .A1(data_in[14]), .A2(n109), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n165), .B2(n99), .A(n128), .ZN(n20) );
  NAND2_X1 U45 ( .A1(data_in[15]), .A2(n109), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n166), .B2(n109), .A(n127), .ZN(n19) );
  NAND2_X1 U47 ( .A1(data_in[16]), .A2(n100), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n167), .B2(n100), .A(n126), .ZN(n18) );
  NAND2_X1 U49 ( .A1(data_in[17]), .A2(n109), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n168), .B2(n109), .A(n125), .ZN(n17) );
  NAND2_X1 U51 ( .A1(data_in[18]), .A2(n99), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n169), .B2(n100), .A(n124), .ZN(n16) );
  NAND2_X1 U53 ( .A1(data_in[19]), .A2(n109), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n170), .B2(n109), .A(n123), .ZN(n15) );
  NAND2_X1 U55 ( .A1(data_in[20]), .A2(n99), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n171), .B2(n99), .A(n122), .ZN(n14) );
  NAND2_X1 U57 ( .A1(data_in[21]), .A2(n109), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n172), .B2(n100), .A(n121), .ZN(n13) );
  NAND2_X1 U59 ( .A1(data_in[22]), .A2(n109), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n173), .B2(n99), .A(n120), .ZN(n12) );
  NAND2_X1 U61 ( .A1(data_in[23]), .A2(n109), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n174), .B2(n99), .A(n119), .ZN(n11) );
  NAND2_X1 U63 ( .A1(data_in[24]), .A2(n100), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n175), .B2(n99), .A(n118), .ZN(n10) );
  NAND2_X1 U65 ( .A1(data_in[25]), .A2(n99), .ZN(n118) );
  CLKBUF_X1 U68 ( .A(rst), .Z(n117) );
  CLKBUF_X1 U70 ( .A(ld), .Z(n99) );
  CLKBUF_X1 U74 ( .A(ld), .Z(n100) );
  CLKBUF_X1 U81 ( .A(ld), .Z(n109) );
  DFFR_X1 \data_out_reg[31]  ( .D(n4), .CK(clk), .RN(n117), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n5), .CK(clk), .RN(n117), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n6), .CK(clk), .RN(n117), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n7), .CK(clk), .RN(n117), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n8), .CK(clk), .RN(n117), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n9), .CK(clk), .RN(n117), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n10), .CK(clk), .RN(n117), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n11), .CK(clk), .RN(n117), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n12), .CK(clk), .RN(n117), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n13), .CK(clk), .RN(n117), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n14), .CK(clk), .RN(n117), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n15), .CK(clk), .RN(n117), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n16), .CK(clk), .RN(n117), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n17), .CK(clk), .RN(n117), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n23), .CK(clk), .RN(n117), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n24), .CK(clk), .RN(n117), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n25), .CK(clk), .RN(rst), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n26), .CK(clk), .RN(rst), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n27), .CK(clk), .RN(rst), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n28), .CK(clk), .RN(rst), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n29), .CK(clk), .RN(rst), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n30), .CK(clk), .RN(rst), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n31), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n33), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n34), .CK(clk), .RN(n117), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n35), .CK(clk), .RN(n117), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N5_0 ( clk, rst, ld, data_in, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  OAI21_X1 U2 ( .B1(n22), .B2(ld), .A(n21), .ZN(n5) );
  NAND2_X1 U3 ( .A1(ld), .A2(data_in[0]), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n23), .B2(ld), .A(n20), .ZN(n4) );
  NAND2_X1 U5 ( .A1(data_in[1]), .A2(ld), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(ld), .A(n19), .ZN(n3) );
  NAND2_X1 U7 ( .A1(data_in[2]), .A2(ld), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n25), .B2(ld), .A(n18), .ZN(n2) );
  NAND2_X1 U9 ( .A1(data_in[3]), .A2(ld), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n26), .B2(ld), .A(n17), .ZN(n1) );
  NAND2_X1 U11 ( .A1(data_in[4]), .A2(ld), .ZN(n17) );
  DFFR_X1 \data_out_reg[4]  ( .D(n1), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n26) );
  DFFR_X1 \data_out_reg[3]  ( .D(n2), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n25) );
  DFFR_X1 \data_out_reg[2]  ( .D(n3), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n24) );
  DFFR_X1 \data_out_reg[1]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n23) );
  DFFR_X1 \data_out_reg[0]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n22) );
endmodule


module reg_file_Dbits32_Abits5 ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n2130, n2135, n2140, n2145, n2150, n2155, n2160, n2165,
         n2170, n2175, n2180, n2185, n2190, n2195, n2200, n2205, n2210, n2215,
         n2220, n2225, n2230, n2235, n2240, n2245, n2250, n2255, n2260, n2265,
         n2270, n2352, n2355, n2358, n2361, n2364, n2367, n2370, n2373, n2376,
         n2379, n2382, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2131, n2132, n2133, n2134, n2136, n2137, n2138,
         n2139, n2141, n2142, n2143, n2144, n2146, n2147, n2148, n2149, n2151,
         n2152, n2153, n2154, n2156, n2157, n2158, n2159, n2161, n2162, n2163,
         n2164, n2166, n2167, n2168, n2169, n2171, n2172, n2173, n2174, n2176,
         n2177, n2178, n2179, n2181, n2182, n2183, n2184, n2186, n2187, n2188,
         n2189, n2191, n2192, n2193, n2194, n2196, n2197, n2198, n2199, n2201,
         n2202, n2203, n2204, n2206, n2207, n2208, n2209, n2211, n2212, n2213,
         n2214, n2216, n2217, n2218, n2219, n2221, n2222, n2223, n2224, n2226,
         n2227, n2228, n2229, n2231, n2232, n2233, n2234, n2236, n2237, n2238,
         n2239, n2241, n2242, n2243, n2244, n2246, n2247, n2248, n2249, n2251,
         n2252, n2253, n2254, n2256, n2257, n2258, n2259, n2261, n2262, n2263,
         n2264, n2266, n2267, n2268, n2269, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2353, n2354, n2356, n2357,
         n2359, n2360, n2362, n2363, n2365, n2366, n2368, n2369, n2371, n2372,
         n2374, n2375, n2377, n2378, n2380, n2381, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5461, n5463,
         n5467, n5470, n5473, n5476, n5477, n5482, n5485, n5488, n5491, n5494,
         n5497, n5500, n5503, n5506, n5507, n5511, n5515, n5518, n5521, n5524,
         n5525, n5530, n5533, n5536, n5539, n5542, n5545, n5547, n5551, n5554,
         n5558, n5560, n5562, n5566, n5570, n5572, n5573, n5578, n5581, n5584,
         n5587, n5590, n5591, n5596, n5598, n5602, n5605, n5608, n5611, n5614,
         n5617, n5620, n5623, n5626, n5629, n5632, n5634, n5638, n5641, n5644,
         n5645, n5650, n5653, n5656, n5659, n5662, n5664, n5668, n5671, n5674,
         n5677, n5680, n5681, n5686, n5689, n5691, n5695, n5698, n5701, n5704,
         n5707, n5709, n5713, n5716, n5717, n5722, n5725, n5728, n5731, n5734,
         n5735, n5740, n5743, n5746, n5749, n5752, n5755, n5758, n5761, n5763,
         n5769, n5770, n5775, n5776, n5781, n5782, n5783, n5785, n5793, n5794,
         n5799, n5800, n5805, n5806, n5807, n5809, n5817, n5818, n5819, n5821,
         n5829, n5830, n5835, n5836, n5840, n5841, n5846, n5847, n5849, n5851,
         n5859, n5860, n5861, n5863, n5868, n5872, n5876, n5877, n5879, n5880,
         n5888, n5889, n5894, n5896, n5898, n5902, n5906, n5907, n5910, n5914,
         n5918, n5920, n5924, n5926, n5928, n5929, n5939, n5946, n5948, n5949,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5974, n5982, n5983, n5984, n5985, n5992, n5993, n6059,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624;

  OAI21_X1 U560 ( .B1(n5928), .B2(n5461), .A(n1488), .ZN(n4189) );
  NAND2_X1 U561 ( .A1(n5929), .A2(n6172), .ZN(n1488) );
  OAI21_X1 U562 ( .B1(n5929), .B2(n6077), .A(n1489), .ZN(n4188) );
  NAND2_X1 U563 ( .A1(n5928), .A2(n6173), .ZN(n1489) );
  OAI21_X1 U564 ( .B1(n5928), .B2(n5467), .A(n1490), .ZN(n4187) );
  NAND2_X1 U565 ( .A1(n5929), .A2(n6174), .ZN(n1490) );
  OAI21_X1 U566 ( .B1(n5929), .B2(n5470), .A(n1491), .ZN(n4186) );
  NAND2_X1 U567 ( .A1(n1487), .A2(n6175), .ZN(n1491) );
  OAI21_X1 U568 ( .B1(n5928), .B2(n5473), .A(n1492), .ZN(n4185) );
  NAND2_X1 U569 ( .A1(n5928), .A2(n6176), .ZN(n1492) );
  OAI21_X1 U570 ( .B1(n5929), .B2(n5476), .A(n1493), .ZN(n4184) );
  NAND2_X1 U571 ( .A1(n1487), .A2(n6177), .ZN(n1493) );
  OAI21_X1 U572 ( .B1(n5928), .B2(n6082), .A(n1494), .ZN(n4183) );
  NAND2_X1 U573 ( .A1(n1487), .A2(n6178), .ZN(n1494) );
  OAI21_X1 U574 ( .B1(n5929), .B2(n5482), .A(n1495), .ZN(n4182) );
  NAND2_X1 U575 ( .A1(n1487), .A2(n6179), .ZN(n1495) );
  OAI21_X1 U576 ( .B1(n5928), .B2(n5485), .A(n1496), .ZN(n4181) );
  NAND2_X1 U577 ( .A1(n1487), .A2(n6180), .ZN(n1496) );
  OAI21_X1 U578 ( .B1(n5929), .B2(n5488), .A(n1497), .ZN(n4180) );
  NAND2_X1 U579 ( .A1(n1487), .A2(n6181), .ZN(n1497) );
  OAI21_X1 U580 ( .B1(n5928), .B2(n5491), .A(n1498), .ZN(n4179) );
  NAND2_X1 U581 ( .A1(n1487), .A2(n6182), .ZN(n1498) );
  OAI21_X1 U582 ( .B1(n5929), .B2(n5494), .A(n1499), .ZN(n4178) );
  NAND2_X1 U583 ( .A1(n1487), .A2(n6183), .ZN(n1499) );
  OAI21_X1 U584 ( .B1(n5928), .B2(n5497), .A(n1500), .ZN(n4177) );
  NAND2_X1 U585 ( .A1(n1487), .A2(n6184), .ZN(n1500) );
  OAI21_X1 U586 ( .B1(n5928), .B2(n5500), .A(n1501), .ZN(n4176) );
  NAND2_X1 U587 ( .A1(n1487), .A2(n6185), .ZN(n1501) );
  OAI21_X1 U588 ( .B1(n5928), .B2(n5503), .A(n1502), .ZN(n4175) );
  NAND2_X1 U589 ( .A1(n1487), .A2(n6186), .ZN(n1502) );
  OAI21_X1 U590 ( .B1(n5928), .B2(n5506), .A(n1503), .ZN(n4174) );
  NAND2_X1 U591 ( .A1(n1487), .A2(n6187), .ZN(n1503) );
  OAI21_X1 U592 ( .B1(n5928), .B2(n6092), .A(n1504), .ZN(n4173) );
  NAND2_X1 U593 ( .A1(n1487), .A2(n6188), .ZN(n1504) );
  OAI21_X1 U594 ( .B1(n5928), .B2(n6093), .A(n1505), .ZN(n4172) );
  NAND2_X1 U595 ( .A1(n5929), .A2(n6189), .ZN(n1505) );
  OAI21_X1 U596 ( .B1(n5928), .B2(n5515), .A(n1506), .ZN(n4171) );
  NAND2_X1 U597 ( .A1(n5928), .A2(n6190), .ZN(n1506) );
  OAI21_X1 U598 ( .B1(n5928), .B2(n5518), .A(n1507), .ZN(n4170) );
  NAND2_X1 U599 ( .A1(n5928), .A2(n6191), .ZN(n1507) );
  OAI21_X1 U600 ( .B1(n5928), .B2(n5521), .A(n1508), .ZN(n4169) );
  NAND2_X1 U601 ( .A1(n5929), .A2(n6192), .ZN(n1508) );
  OAI21_X1 U602 ( .B1(n5928), .B2(n5524), .A(n1509), .ZN(n4168) );
  NAND2_X1 U603 ( .A1(n1487), .A2(n6193), .ZN(n1509) );
  OAI21_X1 U604 ( .B1(n5929), .B2(n6098), .A(n1510), .ZN(n4167) );
  NAND2_X1 U605 ( .A1(n1487), .A2(n6194), .ZN(n1510) );
  OAI21_X1 U606 ( .B1(n5929), .B2(n5530), .A(n1511), .ZN(n4166) );
  NAND2_X1 U607 ( .A1(n1487), .A2(n6195), .ZN(n1511) );
  OAI21_X1 U608 ( .B1(n5929), .B2(n5533), .A(n1512), .ZN(n4165) );
  NAND2_X1 U609 ( .A1(n1487), .A2(n6196), .ZN(n1512) );
  OAI21_X1 U610 ( .B1(n5929), .B2(n5536), .A(n1513), .ZN(n4164) );
  NAND2_X1 U611 ( .A1(n1487), .A2(n6197), .ZN(n1513) );
  OAI21_X1 U612 ( .B1(n5929), .B2(n5539), .A(n1514), .ZN(n4163) );
  NAND2_X1 U613 ( .A1(n1487), .A2(n6198), .ZN(n1514) );
  OAI21_X1 U614 ( .B1(n5929), .B2(n5542), .A(n1515), .ZN(n4162) );
  NAND2_X1 U615 ( .A1(n1487), .A2(n6199), .ZN(n1515) );
  OAI21_X1 U616 ( .B1(n5929), .B2(n5545), .A(n1516), .ZN(n4161) );
  NAND2_X1 U617 ( .A1(n5929), .A2(n6200), .ZN(n1516) );
  OAI21_X1 U618 ( .B1(n5929), .B2(n6105), .A(n1517), .ZN(n4160) );
  NAND2_X1 U619 ( .A1(n1487), .A2(n6201), .ZN(n1517) );
  OAI21_X1 U620 ( .B1(n5929), .B2(n5551), .A(n1518), .ZN(n4159) );
  NAND2_X1 U621 ( .A1(n1487), .A2(n6202), .ZN(n1518) );
  OAI21_X1 U622 ( .B1(n5929), .B2(n5554), .A(n1519), .ZN(n4158) );
  NAND2_X1 U623 ( .A1(n1487), .A2(n6203), .ZN(n1519) );
  NAND2_X1 U624 ( .A1(n1520), .A2(n1521), .ZN(n1487) );
  OAI21_X1 U625 ( .B1(n5461), .B2(n5924), .A(n1523), .ZN(n4157) );
  NAND2_X1 U626 ( .A1(n5924), .A2(n6236), .ZN(n1523) );
  OAI21_X1 U627 ( .B1(n6077), .B2(n5924), .A(n1524), .ZN(n4156) );
  NAND2_X1 U628 ( .A1(n5926), .A2(n6237), .ZN(n1524) );
  OAI21_X1 U629 ( .B1(n5467), .B2(n5924), .A(n1525), .ZN(n4155) );
  NAND2_X1 U630 ( .A1(n5926), .A2(n6238), .ZN(n1525) );
  OAI21_X1 U631 ( .B1(n5470), .B2(n5924), .A(n1526), .ZN(n4154) );
  NAND2_X1 U632 ( .A1(n2270), .A2(n1522), .ZN(n1526) );
  OAI21_X1 U633 ( .B1(n5473), .B2(n5924), .A(n1527), .ZN(n4153) );
  NAND2_X1 U634 ( .A1(n2265), .A2(n1522), .ZN(n1527) );
  OAI21_X1 U635 ( .B1(n5476), .B2(n5924), .A(n1528), .ZN(n4152) );
  NAND2_X1 U636 ( .A1(n2260), .A2(n1522), .ZN(n1528) );
  OAI21_X1 U637 ( .B1(n6082), .B2(n5924), .A(n1529), .ZN(n4151) );
  NAND2_X1 U638 ( .A1(n2255), .A2(n1522), .ZN(n1529) );
  OAI21_X1 U639 ( .B1(n5482), .B2(n5924), .A(n1530), .ZN(n4150) );
  NAND2_X1 U640 ( .A1(n2250), .A2(n5924), .ZN(n1530) );
  OAI21_X1 U641 ( .B1(n5485), .B2(n5924), .A(n1531), .ZN(n4149) );
  NAND2_X1 U642 ( .A1(n2245), .A2(n1522), .ZN(n1531) );
  OAI21_X1 U643 ( .B1(n5488), .B2(n5924), .A(n1532), .ZN(n4148) );
  NAND2_X1 U644 ( .A1(n2240), .A2(n1522), .ZN(n1532) );
  OAI21_X1 U645 ( .B1(n5491), .B2(n5924), .A(n1533), .ZN(n4147) );
  NAND2_X1 U646 ( .A1(n2235), .A2(n1522), .ZN(n1533) );
  OAI21_X1 U647 ( .B1(n5494), .B2(n5924), .A(n1534), .ZN(n4146) );
  NAND2_X1 U648 ( .A1(n2230), .A2(n1522), .ZN(n1534) );
  OAI21_X1 U649 ( .B1(n5497), .B2(n5926), .A(n1535), .ZN(n4145) );
  NAND2_X1 U650 ( .A1(n2225), .A2(n1522), .ZN(n1535) );
  OAI21_X1 U651 ( .B1(n5500), .B2(n5924), .A(n1536), .ZN(n4144) );
  NAND2_X1 U652 ( .A1(n2220), .A2(n5926), .ZN(n1536) );
  OAI21_X1 U653 ( .B1(n5503), .B2(n5926), .A(n1537), .ZN(n4143) );
  NAND2_X1 U654 ( .A1(n2215), .A2(n1522), .ZN(n1537) );
  OAI21_X1 U655 ( .B1(n5506), .B2(n5924), .A(n1538), .ZN(n4142) );
  NAND2_X1 U656 ( .A1(n2210), .A2(n1522), .ZN(n1538) );
  OAI21_X1 U657 ( .B1(n6092), .B2(n5926), .A(n1539), .ZN(n4141) );
  NAND2_X1 U658 ( .A1(n2205), .A2(n5926), .ZN(n1539) );
  OAI21_X1 U659 ( .B1(n6093), .B2(n5924), .A(n1540), .ZN(n4140) );
  NAND2_X1 U660 ( .A1(n2200), .A2(n5924), .ZN(n1540) );
  OAI21_X1 U661 ( .B1(n5515), .B2(n5926), .A(n1541), .ZN(n4139) );
  NAND2_X1 U662 ( .A1(n2195), .A2(n5924), .ZN(n1541) );
  OAI21_X1 U663 ( .B1(n5518), .B2(n5924), .A(n1542), .ZN(n4138) );
  NAND2_X1 U664 ( .A1(n2190), .A2(n1522), .ZN(n1542) );
  OAI21_X1 U665 ( .B1(n5521), .B2(n5926), .A(n1543), .ZN(n4137) );
  NAND2_X1 U666 ( .A1(n2185), .A2(n5926), .ZN(n1543) );
  OAI21_X1 U667 ( .B1(n5524), .B2(n5924), .A(n1544), .ZN(n4136) );
  NAND2_X1 U668 ( .A1(n2180), .A2(n5926), .ZN(n1544) );
  OAI21_X1 U669 ( .B1(n6098), .B2(n5926), .A(n1545), .ZN(n4135) );
  NAND2_X1 U670 ( .A1(n2175), .A2(n1522), .ZN(n1545) );
  OAI21_X1 U671 ( .B1(n5530), .B2(n5926), .A(n1546), .ZN(n4134) );
  NAND2_X1 U672 ( .A1(n2170), .A2(n1522), .ZN(n1546) );
  OAI21_X1 U673 ( .B1(n5533), .B2(n5926), .A(n1547), .ZN(n4133) );
  NAND2_X1 U674 ( .A1(n2165), .A2(n1522), .ZN(n1547) );
  OAI21_X1 U675 ( .B1(n5536), .B2(n5926), .A(n1548), .ZN(n4132) );
  NAND2_X1 U676 ( .A1(n2160), .A2(n1522), .ZN(n1548) );
  OAI21_X1 U677 ( .B1(n5539), .B2(n5926), .A(n1549), .ZN(n4131) );
  NAND2_X1 U678 ( .A1(n2155), .A2(n1522), .ZN(n1549) );
  OAI21_X1 U679 ( .B1(n5542), .B2(n5926), .A(n1550), .ZN(n4130) );
  NAND2_X1 U680 ( .A1(n2150), .A2(n1522), .ZN(n1550) );
  OAI21_X1 U681 ( .B1(n5545), .B2(n5926), .A(n1551), .ZN(n4129) );
  NAND2_X1 U682 ( .A1(n2145), .A2(n1522), .ZN(n1551) );
  OAI21_X1 U683 ( .B1(n6105), .B2(n5926), .A(n1552), .ZN(n4128) );
  NAND2_X1 U684 ( .A1(n2140), .A2(n1522), .ZN(n1552) );
  OAI21_X1 U685 ( .B1(n5551), .B2(n5926), .A(n1553), .ZN(n4127) );
  NAND2_X1 U686 ( .A1(n2135), .A2(n1522), .ZN(n1553) );
  OAI21_X1 U687 ( .B1(n5554), .B2(n5926), .A(n1554), .ZN(n4126) );
  NAND2_X1 U688 ( .A1(n2130), .A2(n1522), .ZN(n1554) );
  NAND2_X1 U689 ( .A1(n1555), .A2(n1556), .ZN(n1522) );
  OAI21_X1 U690 ( .B1(n5461), .B2(n5918), .A(n1558), .ZN(n4125) );
  NAND2_X1 U691 ( .A1(n1557), .A2(n6239), .ZN(n1558) );
  OAI21_X1 U692 ( .B1(n6077), .B2(n5918), .A(n1559), .ZN(n4124) );
  NAND2_X1 U693 ( .A1(n1557), .A2(n6240), .ZN(n1559) );
  OAI21_X1 U694 ( .B1(n5467), .B2(n5918), .A(n1560), .ZN(n4123) );
  NAND2_X1 U695 ( .A1(n1557), .A2(n6241), .ZN(n1560) );
  OAI21_X1 U696 ( .B1(n5470), .B2(n5918), .A(n1561), .ZN(n4122) );
  NAND2_X1 U697 ( .A1(n1557), .A2(n6242), .ZN(n1561) );
  OAI21_X1 U698 ( .B1(n5473), .B2(n5918), .A(n1562), .ZN(n4121) );
  NAND2_X1 U699 ( .A1(n1557), .A2(n6243), .ZN(n1562) );
  OAI21_X1 U700 ( .B1(n5476), .B2(n5918), .A(n1563), .ZN(n4120) );
  NAND2_X1 U701 ( .A1(n1557), .A2(n6244), .ZN(n1563) );
  OAI21_X1 U702 ( .B1(n6082), .B2(n5918), .A(n1564), .ZN(n4119) );
  NAND2_X1 U703 ( .A1(n5920), .A2(n6245), .ZN(n1564) );
  OAI21_X1 U704 ( .B1(n5482), .B2(n5918), .A(n1565), .ZN(n4118) );
  NAND2_X1 U705 ( .A1(n5918), .A2(n6246), .ZN(n1565) );
  OAI21_X1 U706 ( .B1(n5485), .B2(n5918), .A(n1566), .ZN(n4117) );
  NAND2_X1 U707 ( .A1(n5920), .A2(n6247), .ZN(n1566) );
  OAI21_X1 U708 ( .B1(n5488), .B2(n5918), .A(n1567), .ZN(n4116) );
  NAND2_X1 U709 ( .A1(n5918), .A2(n6248), .ZN(n1567) );
  OAI21_X1 U710 ( .B1(n5491), .B2(n5918), .A(n1568), .ZN(n4115) );
  NAND2_X1 U711 ( .A1(n5918), .A2(n6249), .ZN(n1568) );
  OAI21_X1 U712 ( .B1(n5494), .B2(n5918), .A(n1569), .ZN(n4114) );
  NAND2_X1 U713 ( .A1(n1557), .A2(n6250), .ZN(n1569) );
  OAI21_X1 U714 ( .B1(n5497), .B2(n5920), .A(n1570), .ZN(n4113) );
  NAND2_X1 U715 ( .A1(n1557), .A2(n6251), .ZN(n1570) );
  OAI21_X1 U716 ( .B1(n5500), .B2(n5918), .A(n1571), .ZN(n4112) );
  NAND2_X1 U717 ( .A1(n1557), .A2(n6252), .ZN(n1571) );
  OAI21_X1 U718 ( .B1(n5503), .B2(n5920), .A(n1572), .ZN(n4111) );
  NAND2_X1 U719 ( .A1(n1557), .A2(n6253), .ZN(n1572) );
  OAI21_X1 U720 ( .B1(n5506), .B2(n5918), .A(n1573), .ZN(n4110) );
  NAND2_X1 U721 ( .A1(n1557), .A2(n6254), .ZN(n1573) );
  OAI21_X1 U722 ( .B1(n6092), .B2(n5920), .A(n1574), .ZN(n4109) );
  NAND2_X1 U723 ( .A1(n5920), .A2(n6255), .ZN(n1574) );
  OAI21_X1 U724 ( .B1(n6093), .B2(n5918), .A(n1575), .ZN(n4108) );
  NAND2_X1 U725 ( .A1(n1557), .A2(n6256), .ZN(n1575) );
  OAI21_X1 U726 ( .B1(n5515), .B2(n5920), .A(n1576), .ZN(n4107) );
  NAND2_X1 U727 ( .A1(n1557), .A2(n6257), .ZN(n1576) );
  OAI21_X1 U728 ( .B1(n5518), .B2(n5918), .A(n1577), .ZN(n4106) );
  NAND2_X1 U729 ( .A1(n5918), .A2(n6258), .ZN(n1577) );
  OAI21_X1 U730 ( .B1(n5521), .B2(n5920), .A(n1578), .ZN(n4105) );
  NAND2_X1 U731 ( .A1(n5920), .A2(n6259), .ZN(n1578) );
  OAI21_X1 U732 ( .B1(n5524), .B2(n5918), .A(n1579), .ZN(n4104) );
  NAND2_X1 U733 ( .A1(n5920), .A2(n6260), .ZN(n1579) );
  OAI21_X1 U734 ( .B1(n6098), .B2(n5920), .A(n1580), .ZN(n4103) );
  NAND2_X1 U735 ( .A1(n1557), .A2(n6261), .ZN(n1580) );
  OAI21_X1 U736 ( .B1(n5530), .B2(n5920), .A(n1581), .ZN(n4102) );
  NAND2_X1 U737 ( .A1(n1557), .A2(n6262), .ZN(n1581) );
  OAI21_X1 U738 ( .B1(n5533), .B2(n5920), .A(n1582), .ZN(n4101) );
  NAND2_X1 U739 ( .A1(n1557), .A2(n6263), .ZN(n1582) );
  OAI21_X1 U740 ( .B1(n5536), .B2(n5920), .A(n1583), .ZN(n4100) );
  NAND2_X1 U741 ( .A1(n1557), .A2(n6264), .ZN(n1583) );
  OAI21_X1 U742 ( .B1(n5539), .B2(n5920), .A(n1584), .ZN(n4099) );
  NAND2_X1 U743 ( .A1(n1557), .A2(n6265), .ZN(n1584) );
  OAI21_X1 U744 ( .B1(n5542), .B2(n5920), .A(n1585), .ZN(n4098) );
  NAND2_X1 U745 ( .A1(n1557), .A2(n6266), .ZN(n1585) );
  OAI21_X1 U746 ( .B1(n5545), .B2(n5920), .A(n1586), .ZN(n4097) );
  NAND2_X1 U747 ( .A1(n1557), .A2(n6267), .ZN(n1586) );
  OAI21_X1 U748 ( .B1(n6105), .B2(n5920), .A(n1587), .ZN(n4096) );
  NAND2_X1 U749 ( .A1(n1557), .A2(n6268), .ZN(n1587) );
  OAI21_X1 U750 ( .B1(n5551), .B2(n5920), .A(n1588), .ZN(n4095) );
  NAND2_X1 U751 ( .A1(n1557), .A2(n6269), .ZN(n1588) );
  OAI21_X1 U752 ( .B1(n5554), .B2(n5920), .A(n1589), .ZN(n4094) );
  NAND2_X1 U753 ( .A1(n1557), .A2(n6270), .ZN(n1589) );
  NAND2_X1 U754 ( .A1(n1590), .A2(n1556), .ZN(n1557) );
  OAI21_X1 U755 ( .B1(n5461), .B2(n5914), .A(n1592), .ZN(n4093) );
  NAND2_X1 U756 ( .A1(n5914), .A2(n6303), .ZN(n1592) );
  OAI21_X1 U757 ( .B1(n6077), .B2(n5910), .A(n1593), .ZN(n4092) );
  NAND2_X1 U758 ( .A1(n1591), .A2(n6304), .ZN(n1593) );
  OAI21_X1 U759 ( .B1(n5467), .B2(n5914), .A(n1594), .ZN(n4091) );
  NAND2_X1 U760 ( .A1(n5910), .A2(n6305), .ZN(n1594) );
  OAI21_X1 U761 ( .B1(n5470), .B2(n5910), .A(n1595), .ZN(n4090) );
  NAND2_X1 U762 ( .A1(n5914), .A2(n6306), .ZN(n1595) );
  OAI21_X1 U763 ( .B1(n5473), .B2(n5914), .A(n1596), .ZN(n4089) );
  NAND2_X1 U764 ( .A1(n5910), .A2(n6307), .ZN(n1596) );
  OAI21_X1 U765 ( .B1(n5476), .B2(n5910), .A(n1597), .ZN(n4088) );
  NAND2_X1 U766 ( .A1(n5910), .A2(n6308), .ZN(n1597) );
  OAI21_X1 U767 ( .B1(n6082), .B2(n5914), .A(n1598), .ZN(n4087) );
  NAND2_X1 U768 ( .A1(n5910), .A2(n6309), .ZN(n1598) );
  OAI21_X1 U769 ( .B1(n5482), .B2(n5910), .A(n1599), .ZN(n4086) );
  NAND2_X1 U770 ( .A1(n1591), .A2(n6310), .ZN(n1599) );
  OAI21_X1 U771 ( .B1(n5485), .B2(n5914), .A(n1600), .ZN(n4085) );
  NAND2_X1 U772 ( .A1(n1591), .A2(n6311), .ZN(n1600) );
  OAI21_X1 U773 ( .B1(n5488), .B2(n5910), .A(n1601), .ZN(n4084) );
  NAND2_X1 U774 ( .A1(n1591), .A2(n6312), .ZN(n1601) );
  OAI21_X1 U775 ( .B1(n5491), .B2(n5914), .A(n1602), .ZN(n4083) );
  NAND2_X1 U776 ( .A1(n1591), .A2(n6313), .ZN(n1602) );
  OAI21_X1 U777 ( .B1(n5494), .B2(n5914), .A(n1603), .ZN(n4082) );
  NAND2_X1 U778 ( .A1(n1591), .A2(n6314), .ZN(n1603) );
  OAI21_X1 U779 ( .B1(n5497), .B2(n5910), .A(n1604), .ZN(n4081) );
  NAND2_X1 U780 ( .A1(n1591), .A2(n6315), .ZN(n1604) );
  OAI21_X1 U781 ( .B1(n5500), .B2(n5910), .A(n1605), .ZN(n4080) );
  NAND2_X1 U782 ( .A1(n1591), .A2(n6316), .ZN(n1605) );
  OAI21_X1 U783 ( .B1(n5503), .B2(n5914), .A(n1606), .ZN(n4079) );
  NAND2_X1 U784 ( .A1(n1591), .A2(n6317), .ZN(n1606) );
  OAI21_X1 U785 ( .B1(n5506), .B2(n5910), .A(n1607), .ZN(n4078) );
  NAND2_X1 U786 ( .A1(n1591), .A2(n6318), .ZN(n1607) );
  OAI21_X1 U787 ( .B1(n6092), .B2(n1591), .A(n1608), .ZN(n4077) );
  NAND2_X1 U788 ( .A1(n5910), .A2(n6319), .ZN(n1608) );
  OAI21_X1 U789 ( .B1(n6093), .B2(n1591), .A(n1609), .ZN(n4076) );
  NAND2_X1 U790 ( .A1(n1591), .A2(n6320), .ZN(n1609) );
  OAI21_X1 U791 ( .B1(n5515), .B2(n1591), .A(n1610), .ZN(n4075) );
  NAND2_X1 U792 ( .A1(n5910), .A2(n6321), .ZN(n1610) );
  OAI21_X1 U793 ( .B1(n5518), .B2(n1591), .A(n1611), .ZN(n4074) );
  NAND2_X1 U794 ( .A1(n5910), .A2(n6322), .ZN(n1611) );
  OAI21_X1 U795 ( .B1(n5521), .B2(n1591), .A(n1612), .ZN(n4073) );
  NAND2_X1 U796 ( .A1(n5910), .A2(n6323), .ZN(n1612) );
  OAI21_X1 U797 ( .B1(n5524), .B2(n1591), .A(n1613), .ZN(n4072) );
  NAND2_X1 U798 ( .A1(n5910), .A2(n6324), .ZN(n1613) );
  OAI21_X1 U799 ( .B1(n6098), .B2(n5914), .A(n1614), .ZN(n4071) );
  NAND2_X1 U800 ( .A1(n5910), .A2(n6325), .ZN(n1614) );
  OAI21_X1 U801 ( .B1(n5530), .B2(n5914), .A(n1615), .ZN(n4070) );
  NAND2_X1 U802 ( .A1(n5910), .A2(n6326), .ZN(n1615) );
  OAI21_X1 U803 ( .B1(n5533), .B2(n5914), .A(n1616), .ZN(n4069) );
  NAND2_X1 U804 ( .A1(n5910), .A2(n6327), .ZN(n1616) );
  OAI21_X1 U805 ( .B1(n5536), .B2(n5914), .A(n1617), .ZN(n4068) );
  NAND2_X1 U806 ( .A1(n1591), .A2(n6328), .ZN(n1617) );
  OAI21_X1 U807 ( .B1(n5539), .B2(n5914), .A(n1618), .ZN(n4067) );
  NAND2_X1 U808 ( .A1(n1591), .A2(n6329), .ZN(n1618) );
  OAI21_X1 U809 ( .B1(n5542), .B2(n5914), .A(n1619), .ZN(n4066) );
  NAND2_X1 U810 ( .A1(n1591), .A2(n6330), .ZN(n1619) );
  OAI21_X1 U811 ( .B1(n5545), .B2(n5914), .A(n1620), .ZN(n4065) );
  NAND2_X1 U812 ( .A1(n1591), .A2(n6331), .ZN(n1620) );
  OAI21_X1 U813 ( .B1(n6105), .B2(n5914), .A(n1621), .ZN(n4064) );
  NAND2_X1 U814 ( .A1(n5910), .A2(n6332), .ZN(n1621) );
  OAI21_X1 U815 ( .B1(n5551), .B2(n5914), .A(n1622), .ZN(n4063) );
  NAND2_X1 U816 ( .A1(n1591), .A2(n6333), .ZN(n1622) );
  OAI21_X1 U817 ( .B1(n5554), .B2(n1591), .A(n1623), .ZN(n4062) );
  NAND2_X1 U818 ( .A1(n5914), .A2(n6334), .ZN(n1623) );
  NAND2_X1 U819 ( .A1(n1624), .A2(n1556), .ZN(n1591) );
  OAI21_X1 U820 ( .B1(n5461), .B2(n5906), .A(n1626), .ZN(n4061) );
  NAND2_X1 U821 ( .A1(n2382), .A2(n1625), .ZN(n1626) );
  OAI21_X1 U822 ( .B1(n6077), .B2(n5906), .A(n1627), .ZN(n4060) );
  NAND2_X1 U823 ( .A1(n2379), .A2(n1625), .ZN(n1627) );
  OAI21_X1 U824 ( .B1(n5467), .B2(n5906), .A(n1628), .ZN(n4059) );
  NAND2_X1 U825 ( .A1(n2376), .A2(n1625), .ZN(n1628) );
  OAI21_X1 U826 ( .B1(n5470), .B2(n5906), .A(n1629), .ZN(n4058) );
  NAND2_X1 U827 ( .A1(n2373), .A2(n1625), .ZN(n1629) );
  OAI21_X1 U828 ( .B1(n5473), .B2(n5906), .A(n1630), .ZN(n4057) );
  NAND2_X1 U829 ( .A1(n2370), .A2(n1625), .ZN(n1630) );
  OAI21_X1 U830 ( .B1(n5476), .B2(n5906), .A(n1631), .ZN(n4056) );
  NAND2_X1 U831 ( .A1(n2367), .A2(n1625), .ZN(n1631) );
  OAI21_X1 U832 ( .B1(n6082), .B2(n5906), .A(n1632), .ZN(n4055) );
  NAND2_X1 U833 ( .A1(n2364), .A2(n1625), .ZN(n1632) );
  OAI21_X1 U834 ( .B1(n5482), .B2(n5906), .A(n1633), .ZN(n4054) );
  NAND2_X1 U835 ( .A1(n2361), .A2(n1625), .ZN(n1633) );
  OAI21_X1 U836 ( .B1(n5485), .B2(n5906), .A(n1634), .ZN(n4053) );
  NAND2_X1 U837 ( .A1(n2358), .A2(n1625), .ZN(n1634) );
  OAI21_X1 U838 ( .B1(n5488), .B2(n5906), .A(n1635), .ZN(n4052) );
  NAND2_X1 U839 ( .A1(n2355), .A2(n1625), .ZN(n1635) );
  OAI21_X1 U840 ( .B1(n5491), .B2(n5906), .A(n1636), .ZN(n4051) );
  NAND2_X1 U841 ( .A1(n2352), .A2(n1625), .ZN(n1636) );
  OAI21_X1 U842 ( .B1(n5494), .B2(n5907), .A(n1637), .ZN(n4050) );
  NAND2_X1 U843 ( .A1(n5907), .A2(n6335), .ZN(n1637) );
  OAI21_X1 U844 ( .B1(n5497), .B2(n5907), .A(n1638), .ZN(n4049) );
  NAND2_X1 U845 ( .A1(n5906), .A2(n6336), .ZN(n1638) );
  OAI21_X1 U846 ( .B1(n5500), .B2(n5907), .A(n1639), .ZN(n4048) );
  NAND2_X1 U847 ( .A1(n5907), .A2(n6337), .ZN(n1639) );
  OAI21_X1 U848 ( .B1(n5503), .B2(n5907), .A(n1640), .ZN(n4047) );
  NAND2_X1 U849 ( .A1(n5906), .A2(n6338), .ZN(n1640) );
  OAI21_X1 U850 ( .B1(n5506), .B2(n5907), .A(n1641), .ZN(n4046) );
  NAND2_X1 U851 ( .A1(n5907), .A2(n6339), .ZN(n1641) );
  OAI21_X1 U852 ( .B1(n6092), .B2(n5907), .A(n1642), .ZN(n4045) );
  NAND2_X1 U853 ( .A1(n5906), .A2(n6340), .ZN(n1642) );
  OAI21_X1 U854 ( .B1(n6093), .B2(n5907), .A(n1643), .ZN(n4044) );
  NAND2_X1 U855 ( .A1(n5907), .A2(n6341), .ZN(n1643) );
  OAI21_X1 U856 ( .B1(n5515), .B2(n5907), .A(n1644), .ZN(n4043) );
  NAND2_X1 U857 ( .A1(n5906), .A2(n6342), .ZN(n1644) );
  OAI21_X1 U858 ( .B1(n5518), .B2(n5907), .A(n1645), .ZN(n4042) );
  NAND2_X1 U859 ( .A1(n1625), .A2(n6343), .ZN(n1645) );
  OAI21_X1 U860 ( .B1(n5521), .B2(n5907), .A(n1646), .ZN(n4041) );
  NAND2_X1 U861 ( .A1(n1625), .A2(n6344), .ZN(n1646) );
  OAI21_X1 U862 ( .B1(n5524), .B2(n5907), .A(n1647), .ZN(n4040) );
  NAND2_X1 U863 ( .A1(n1625), .A2(n6345), .ZN(n1647) );
  OAI21_X1 U864 ( .B1(n6098), .B2(n5907), .A(n1648), .ZN(n4039) );
  NAND2_X1 U865 ( .A1(n1625), .A2(n6346), .ZN(n1648) );
  OAI21_X1 U866 ( .B1(n5530), .B2(n5907), .A(n1649), .ZN(n4038) );
  NAND2_X1 U867 ( .A1(n1625), .A2(n6347), .ZN(n1649) );
  OAI21_X1 U868 ( .B1(n5533), .B2(n5906), .A(n1650), .ZN(n4037) );
  NAND2_X1 U869 ( .A1(n1625), .A2(n6348), .ZN(n1650) );
  OAI21_X1 U870 ( .B1(n5536), .B2(n5907), .A(n1651), .ZN(n4036) );
  NAND2_X1 U871 ( .A1(n1625), .A2(n6349), .ZN(n1651) );
  OAI21_X1 U872 ( .B1(n5539), .B2(n5906), .A(n1652), .ZN(n4035) );
  NAND2_X1 U873 ( .A1(n1625), .A2(n6350), .ZN(n1652) );
  OAI21_X1 U874 ( .B1(n5542), .B2(n5907), .A(n1653), .ZN(n4034) );
  NAND2_X1 U875 ( .A1(n1625), .A2(n6351), .ZN(n1653) );
  OAI21_X1 U876 ( .B1(n5545), .B2(n5906), .A(n1654), .ZN(n4033) );
  NAND2_X1 U877 ( .A1(n1625), .A2(n6352), .ZN(n1654) );
  OAI21_X1 U878 ( .B1(n6105), .B2(n5907), .A(n1655), .ZN(n4032) );
  NAND2_X1 U879 ( .A1(n5906), .A2(n6353), .ZN(n1655) );
  OAI21_X1 U880 ( .B1(n5551), .B2(n5906), .A(n1656), .ZN(n4031) );
  NAND2_X1 U881 ( .A1(n1625), .A2(n6354), .ZN(n1656) );
  OAI21_X1 U882 ( .B1(n5554), .B2(n5907), .A(n1657), .ZN(n4030) );
  NAND2_X1 U883 ( .A1(n1625), .A2(n6355), .ZN(n1657) );
  NAND2_X1 U884 ( .A1(n1658), .A2(n1556), .ZN(n1625) );
  OAI21_X1 U885 ( .B1(n5461), .B2(n5902), .A(n1660), .ZN(n4029) );
  NAND2_X1 U886 ( .A1(n5902), .A2(n6388), .ZN(n1660) );
  OAI21_X1 U887 ( .B1(n6077), .B2(n5898), .A(n1661), .ZN(n4028) );
  NAND2_X1 U888 ( .A1(n1659), .A2(n6389), .ZN(n1661) );
  OAI21_X1 U889 ( .B1(n5467), .B2(n5902), .A(n1662), .ZN(n4027) );
  NAND2_X1 U890 ( .A1(n5898), .A2(n6390), .ZN(n1662) );
  OAI21_X1 U891 ( .B1(n5470), .B2(n5898), .A(n1663), .ZN(n4026) );
  NAND2_X1 U892 ( .A1(n5902), .A2(n6391), .ZN(n1663) );
  OAI21_X1 U893 ( .B1(n5473), .B2(n5902), .A(n1664), .ZN(n4025) );
  NAND2_X1 U894 ( .A1(n5898), .A2(n6392), .ZN(n1664) );
  OAI21_X1 U895 ( .B1(n5476), .B2(n5898), .A(n1665), .ZN(n4024) );
  NAND2_X1 U896 ( .A1(n5898), .A2(n6393), .ZN(n1665) );
  OAI21_X1 U897 ( .B1(n6082), .B2(n5902), .A(n1666), .ZN(n4023) );
  NAND2_X1 U898 ( .A1(n5898), .A2(n6394), .ZN(n1666) );
  OAI21_X1 U899 ( .B1(n5482), .B2(n5898), .A(n1667), .ZN(n4022) );
  NAND2_X1 U900 ( .A1(n1659), .A2(n6395), .ZN(n1667) );
  OAI21_X1 U901 ( .B1(n5485), .B2(n5902), .A(n1668), .ZN(n4021) );
  NAND2_X1 U902 ( .A1(n1659), .A2(n6396), .ZN(n1668) );
  OAI21_X1 U903 ( .B1(n5488), .B2(n5898), .A(n1669), .ZN(n4020) );
  NAND2_X1 U904 ( .A1(n1659), .A2(n6397), .ZN(n1669) );
  OAI21_X1 U905 ( .B1(n5491), .B2(n5902), .A(n1670), .ZN(n4019) );
  NAND2_X1 U906 ( .A1(n1659), .A2(n6398), .ZN(n1670) );
  OAI21_X1 U907 ( .B1(n5494), .B2(n5902), .A(n1671), .ZN(n4018) );
  NAND2_X1 U908 ( .A1(n1659), .A2(n6399), .ZN(n1671) );
  OAI21_X1 U909 ( .B1(n5497), .B2(n5898), .A(n1672), .ZN(n4017) );
  NAND2_X1 U910 ( .A1(n1659), .A2(n6400), .ZN(n1672) );
  OAI21_X1 U911 ( .B1(n5500), .B2(n5898), .A(n1673), .ZN(n4016) );
  NAND2_X1 U912 ( .A1(n1659), .A2(n6401), .ZN(n1673) );
  OAI21_X1 U913 ( .B1(n5503), .B2(n5902), .A(n1674), .ZN(n4015) );
  NAND2_X1 U914 ( .A1(n1659), .A2(n6402), .ZN(n1674) );
  OAI21_X1 U915 ( .B1(n5506), .B2(n5898), .A(n1675), .ZN(n4014) );
  NAND2_X1 U916 ( .A1(n1659), .A2(n6403), .ZN(n1675) );
  OAI21_X1 U917 ( .B1(n6092), .B2(n1659), .A(n1676), .ZN(n4013) );
  NAND2_X1 U918 ( .A1(n5898), .A2(n6404), .ZN(n1676) );
  OAI21_X1 U919 ( .B1(n6093), .B2(n1659), .A(n1677), .ZN(n4012) );
  NAND2_X1 U920 ( .A1(n1659), .A2(n6405), .ZN(n1677) );
  OAI21_X1 U921 ( .B1(n5515), .B2(n1659), .A(n1678), .ZN(n4011) );
  NAND2_X1 U922 ( .A1(n5898), .A2(n6406), .ZN(n1678) );
  OAI21_X1 U923 ( .B1(n5518), .B2(n1659), .A(n1679), .ZN(n4010) );
  NAND2_X1 U924 ( .A1(n5898), .A2(n6407), .ZN(n1679) );
  OAI21_X1 U925 ( .B1(n5521), .B2(n1659), .A(n1680), .ZN(n4009) );
  NAND2_X1 U926 ( .A1(n5898), .A2(n6408), .ZN(n1680) );
  OAI21_X1 U927 ( .B1(n5524), .B2(n1659), .A(n1681), .ZN(n4008) );
  NAND2_X1 U928 ( .A1(n5898), .A2(n6409), .ZN(n1681) );
  OAI21_X1 U929 ( .B1(n6098), .B2(n5902), .A(n1682), .ZN(n4007) );
  NAND2_X1 U930 ( .A1(n5898), .A2(n6410), .ZN(n1682) );
  OAI21_X1 U931 ( .B1(n5530), .B2(n5902), .A(n1683), .ZN(n4006) );
  NAND2_X1 U932 ( .A1(n5898), .A2(n6411), .ZN(n1683) );
  OAI21_X1 U933 ( .B1(n5533), .B2(n5902), .A(n1684), .ZN(n4005) );
  NAND2_X1 U934 ( .A1(n5898), .A2(n6412), .ZN(n1684) );
  OAI21_X1 U935 ( .B1(n5536), .B2(n5902), .A(n1685), .ZN(n4004) );
  NAND2_X1 U936 ( .A1(n1659), .A2(n6413), .ZN(n1685) );
  OAI21_X1 U937 ( .B1(n5539), .B2(n5902), .A(n1686), .ZN(n4003) );
  NAND2_X1 U938 ( .A1(n1659), .A2(n6414), .ZN(n1686) );
  OAI21_X1 U939 ( .B1(n5542), .B2(n5902), .A(n1687), .ZN(n4002) );
  NAND2_X1 U940 ( .A1(n1659), .A2(n6415), .ZN(n1687) );
  OAI21_X1 U941 ( .B1(n5545), .B2(n5902), .A(n1688), .ZN(n4001) );
  NAND2_X1 U942 ( .A1(n1659), .A2(n6416), .ZN(n1688) );
  OAI21_X1 U943 ( .B1(n6105), .B2(n5902), .A(n1689), .ZN(n4000) );
  NAND2_X1 U944 ( .A1(n5898), .A2(n6417), .ZN(n1689) );
  OAI21_X1 U945 ( .B1(n5551), .B2(n5902), .A(n1690), .ZN(n3999) );
  NAND2_X1 U946 ( .A1(n1659), .A2(n6418), .ZN(n1690) );
  OAI21_X1 U947 ( .B1(n5554), .B2(n1659), .A(n1691), .ZN(n3998) );
  NAND2_X1 U948 ( .A1(n5902), .A2(n6419), .ZN(n1691) );
  NAND2_X1 U949 ( .A1(n1692), .A2(n1555), .ZN(n1659) );
  OAI21_X1 U950 ( .B1(n5461), .B2(n5894), .A(n1694), .ZN(n3918) );
  NAND2_X1 U951 ( .A1(n1693), .A2(n6484), .ZN(n1694) );
  OAI21_X1 U952 ( .B1(n6077), .B2(n5894), .A(n1695), .ZN(n3917) );
  NAND2_X1 U953 ( .A1(n1693), .A2(n6485), .ZN(n1695) );
  OAI21_X1 U954 ( .B1(n5467), .B2(n5894), .A(n1696), .ZN(n3916) );
  NAND2_X1 U955 ( .A1(n1693), .A2(n6486), .ZN(n1696) );
  OAI21_X1 U956 ( .B1(n5470), .B2(n5894), .A(n1697), .ZN(n3915) );
  NAND2_X1 U957 ( .A1(n1693), .A2(n6487), .ZN(n1697) );
  OAI21_X1 U958 ( .B1(n5473), .B2(n5894), .A(n1698), .ZN(n3914) );
  NAND2_X1 U959 ( .A1(n1693), .A2(n6488), .ZN(n1698) );
  OAI21_X1 U960 ( .B1(n5476), .B2(n5894), .A(n1699), .ZN(n3913) );
  NAND2_X1 U961 ( .A1(n1693), .A2(n6489), .ZN(n1699) );
  OAI21_X1 U962 ( .B1(n6082), .B2(n5894), .A(n1700), .ZN(n3912) );
  NAND2_X1 U963 ( .A1(n5896), .A2(n6490), .ZN(n1700) );
  OAI21_X1 U964 ( .B1(n5482), .B2(n5894), .A(n1701), .ZN(n3911) );
  NAND2_X1 U965 ( .A1(n5894), .A2(n6491), .ZN(n1701) );
  OAI21_X1 U966 ( .B1(n5485), .B2(n5894), .A(n1702), .ZN(n3910) );
  NAND2_X1 U967 ( .A1(n5896), .A2(n6492), .ZN(n1702) );
  OAI21_X1 U968 ( .B1(n5488), .B2(n5894), .A(n1703), .ZN(n3909) );
  NAND2_X1 U969 ( .A1(n5894), .A2(n6493), .ZN(n1703) );
  OAI21_X1 U970 ( .B1(n5491), .B2(n5894), .A(n1704), .ZN(n3908) );
  NAND2_X1 U971 ( .A1(n5894), .A2(n6494), .ZN(n1704) );
  OAI21_X1 U972 ( .B1(n5494), .B2(n5894), .A(n1705), .ZN(n3907) );
  NAND2_X1 U973 ( .A1(n1693), .A2(n6495), .ZN(n1705) );
  OAI21_X1 U974 ( .B1(n5497), .B2(n5896), .A(n1706), .ZN(n3906) );
  NAND2_X1 U975 ( .A1(n1693), .A2(n6496), .ZN(n1706) );
  OAI21_X1 U976 ( .B1(n5500), .B2(n5894), .A(n1707), .ZN(n3905) );
  NAND2_X1 U977 ( .A1(n1693), .A2(n6497), .ZN(n1707) );
  OAI21_X1 U978 ( .B1(n5503), .B2(n5896), .A(n1708), .ZN(n3904) );
  NAND2_X1 U979 ( .A1(n1693), .A2(n6498), .ZN(n1708) );
  OAI21_X1 U980 ( .B1(n5506), .B2(n5894), .A(n1709), .ZN(n3903) );
  NAND2_X1 U981 ( .A1(n1693), .A2(n6499), .ZN(n1709) );
  OAI21_X1 U982 ( .B1(n6092), .B2(n5896), .A(n1710), .ZN(n3902) );
  NAND2_X1 U983 ( .A1(n5896), .A2(n6500), .ZN(n1710) );
  OAI21_X1 U984 ( .B1(n6093), .B2(n5894), .A(n1711), .ZN(n3901) );
  NAND2_X1 U985 ( .A1(n1693), .A2(n6501), .ZN(n1711) );
  OAI21_X1 U986 ( .B1(n5515), .B2(n5896), .A(n1712), .ZN(n3900) );
  NAND2_X1 U987 ( .A1(n1693), .A2(n6502), .ZN(n1712) );
  OAI21_X1 U988 ( .B1(n5518), .B2(n5894), .A(n1713), .ZN(n3899) );
  NAND2_X1 U989 ( .A1(n5894), .A2(n6503), .ZN(n1713) );
  OAI21_X1 U990 ( .B1(n5521), .B2(n5896), .A(n1714), .ZN(n3898) );
  NAND2_X1 U991 ( .A1(n5896), .A2(n6504), .ZN(n1714) );
  OAI21_X1 U992 ( .B1(n5524), .B2(n5894), .A(n1715), .ZN(n3897) );
  NAND2_X1 U993 ( .A1(n5896), .A2(n6505), .ZN(n1715) );
  OAI21_X1 U994 ( .B1(n6098), .B2(n5896), .A(n1716), .ZN(n3896) );
  NAND2_X1 U995 ( .A1(n1693), .A2(n6506), .ZN(n1716) );
  OAI21_X1 U996 ( .B1(n5530), .B2(n5896), .A(n1717), .ZN(n3895) );
  NAND2_X1 U997 ( .A1(n1693), .A2(n6507), .ZN(n1717) );
  OAI21_X1 U998 ( .B1(n5533), .B2(n5896), .A(n1718), .ZN(n3894) );
  NAND2_X1 U999 ( .A1(n1693), .A2(n6508), .ZN(n1718) );
  OAI21_X1 U1000 ( .B1(n5536), .B2(n5896), .A(n1719), .ZN(n3893) );
  NAND2_X1 U1001 ( .A1(n1693), .A2(n6509), .ZN(n1719) );
  OAI21_X1 U1002 ( .B1(n5539), .B2(n5896), .A(n1720), .ZN(n3892) );
  NAND2_X1 U1003 ( .A1(n1693), .A2(n6510), .ZN(n1720) );
  OAI21_X1 U1004 ( .B1(n5542), .B2(n5896), .A(n1721), .ZN(n3891) );
  NAND2_X1 U1005 ( .A1(n1693), .A2(n6511), .ZN(n1721) );
  OAI21_X1 U1006 ( .B1(n5545), .B2(n5896), .A(n1722), .ZN(n3890) );
  NAND2_X1 U1007 ( .A1(n1693), .A2(n6512), .ZN(n1722) );
  OAI21_X1 U1008 ( .B1(n6105), .B2(n5896), .A(n1723), .ZN(n3889) );
  NAND2_X1 U1009 ( .A1(n1693), .A2(n6513), .ZN(n1723) );
  OAI21_X1 U1010 ( .B1(n5551), .B2(n5896), .A(n1724), .ZN(n3888) );
  NAND2_X1 U1011 ( .A1(n1693), .A2(n6514), .ZN(n1724) );
  OAI21_X1 U1012 ( .B1(n5554), .B2(n5896), .A(n1725), .ZN(n3887) );
  NAND2_X1 U1013 ( .A1(n1693), .A2(n6515), .ZN(n1725) );
  NAND2_X1 U1014 ( .A1(n1692), .A2(n1658), .ZN(n1693) );
  OAI21_X1 U1015 ( .B1(n5461), .B2(n5888), .A(n1727), .ZN(n3886) );
  NAND2_X1 U1016 ( .A1(n1726), .A2(n6452), .ZN(n1727) );
  OAI21_X1 U1017 ( .B1(n6077), .B2(n5888), .A(n1728), .ZN(n3885) );
  NAND2_X1 U1018 ( .A1(n1726), .A2(n6453), .ZN(n1728) );
  OAI21_X1 U1019 ( .B1(n5467), .B2(n5888), .A(n1729), .ZN(n3884) );
  NAND2_X1 U1020 ( .A1(n1726), .A2(n6454), .ZN(n1729) );
  OAI21_X1 U1021 ( .B1(n5470), .B2(n5888), .A(n1730), .ZN(n3883) );
  NAND2_X1 U1022 ( .A1(n1726), .A2(n6455), .ZN(n1730) );
  OAI21_X1 U1023 ( .B1(n5473), .B2(n5888), .A(n1731), .ZN(n3882) );
  NAND2_X1 U1024 ( .A1(n1726), .A2(n6456), .ZN(n1731) );
  OAI21_X1 U1025 ( .B1(n5476), .B2(n5888), .A(n1732), .ZN(n3881) );
  NAND2_X1 U1026 ( .A1(n1726), .A2(n6457), .ZN(n1732) );
  OAI21_X1 U1027 ( .B1(n6082), .B2(n5888), .A(n1733), .ZN(n3880) );
  NAND2_X1 U1028 ( .A1(n1726), .A2(n6458), .ZN(n1733) );
  OAI21_X1 U1029 ( .B1(n5482), .B2(n5888), .A(n1734), .ZN(n3879) );
  NAND2_X1 U1030 ( .A1(n5889), .A2(n6459), .ZN(n1734) );
  OAI21_X1 U1031 ( .B1(n5485), .B2(n5888), .A(n1735), .ZN(n3878) );
  NAND2_X1 U1032 ( .A1(n5888), .A2(n6460), .ZN(n1735) );
  OAI21_X1 U1033 ( .B1(n5488), .B2(n5888), .A(n1736), .ZN(n3877) );
  NAND2_X1 U1034 ( .A1(n5889), .A2(n6461), .ZN(n1736) );
  OAI21_X1 U1035 ( .B1(n5491), .B2(n5888), .A(n1737), .ZN(n3876) );
  NAND2_X1 U1036 ( .A1(n5888), .A2(n6462), .ZN(n1737) );
  OAI21_X1 U1037 ( .B1(n5494), .B2(n5889), .A(n1738), .ZN(n3875) );
  NAND2_X1 U1038 ( .A1(n5889), .A2(n6463), .ZN(n1738) );
  OAI21_X1 U1039 ( .B1(n5497), .B2(n5889), .A(n1739), .ZN(n3874) );
  NAND2_X1 U1040 ( .A1(n5888), .A2(n6464), .ZN(n1739) );
  OAI21_X1 U1041 ( .B1(n5500), .B2(n5889), .A(n1740), .ZN(n3873) );
  NAND2_X1 U1042 ( .A1(n5889), .A2(n6465), .ZN(n1740) );
  OAI21_X1 U1043 ( .B1(n5503), .B2(n5889), .A(n1741), .ZN(n3872) );
  NAND2_X1 U1044 ( .A1(n5888), .A2(n6466), .ZN(n1741) );
  OAI21_X1 U1045 ( .B1(n5506), .B2(n5889), .A(n1742), .ZN(n3871) );
  NAND2_X1 U1046 ( .A1(n1726), .A2(n6467), .ZN(n1742) );
  OAI21_X1 U1047 ( .B1(n6092), .B2(n5889), .A(n1743), .ZN(n3870) );
  NAND2_X1 U1048 ( .A1(n1726), .A2(n6468), .ZN(n1743) );
  OAI21_X1 U1049 ( .B1(n5461), .B2(n5879), .A(n1745), .ZN(n3869) );
  NAND2_X1 U1050 ( .A1(n2830), .A2(n5879), .ZN(n1745) );
  OAI21_X1 U1051 ( .B1(n6077), .B2(n5880), .A(n1746), .ZN(n3868) );
  NAND2_X1 U1052 ( .A1(n2829), .A2(n5879), .ZN(n1746) );
  OAI21_X1 U1053 ( .B1(n5467), .B2(n1744), .A(n1747), .ZN(n3867) );
  NAND2_X1 U1054 ( .A1(n2828), .A2(n5879), .ZN(n1747) );
  OAI21_X1 U1055 ( .B1(n5470), .B2(n1744), .A(n1748), .ZN(n3866) );
  NAND2_X1 U1056 ( .A1(n2827), .A2(n5879), .ZN(n1748) );
  OAI21_X1 U1057 ( .B1(n5473), .B2(n1744), .A(n1749), .ZN(n3865) );
  NAND2_X1 U1058 ( .A1(n2826), .A2(n5880), .ZN(n1749) );
  OAI21_X1 U1059 ( .B1(n5476), .B2(n1744), .A(n1750), .ZN(n3864) );
  NAND2_X1 U1060 ( .A1(n2825), .A2(n5879), .ZN(n1750) );
  OAI21_X1 U1061 ( .B1(n6082), .B2(n1744), .A(n1751), .ZN(n3863) );
  NAND2_X1 U1062 ( .A1(n2824), .A2(n5879), .ZN(n1751) );
  OAI21_X1 U1063 ( .B1(n5482), .B2(n1744), .A(n1752), .ZN(n3862) );
  NAND2_X1 U1064 ( .A1(n2823), .A2(n5880), .ZN(n1752) );
  OAI21_X1 U1065 ( .B1(n5485), .B2(n1744), .A(n1753), .ZN(n3861) );
  NAND2_X1 U1066 ( .A1(n2822), .A2(n5880), .ZN(n1753) );
  OAI21_X1 U1067 ( .B1(n5488), .B2(n1744), .A(n1754), .ZN(n3860) );
  NAND2_X1 U1068 ( .A1(n2821), .A2(n5880), .ZN(n1754) );
  OAI21_X1 U1069 ( .B1(n5491), .B2(n1744), .A(n1755), .ZN(n3859) );
  NAND2_X1 U1070 ( .A1(n2820), .A2(n5880), .ZN(n1755) );
  OAI21_X1 U1071 ( .B1(n5494), .B2(n1744), .A(n1756), .ZN(n3858) );
  NAND2_X1 U1072 ( .A1(n2819), .A2(n5879), .ZN(n1756) );
  OAI21_X1 U1073 ( .B1(n5497), .B2(n1744), .A(n1757), .ZN(n3857) );
  NAND2_X1 U1074 ( .A1(n2818), .A2(n1744), .ZN(n1757) );
  OAI21_X1 U1075 ( .B1(n5500), .B2(n1744), .A(n1758), .ZN(n3856) );
  NAND2_X1 U1076 ( .A1(n2817), .A2(n5880), .ZN(n1758) );
  OAI21_X1 U1077 ( .B1(n5503), .B2(n1744), .A(n1759), .ZN(n3855) );
  NAND2_X1 U1078 ( .A1(n2816), .A2(n5879), .ZN(n1759) );
  OAI21_X1 U1079 ( .B1(n5506), .B2(n1744), .A(n1760), .ZN(n3854) );
  NAND2_X1 U1080 ( .A1(n2815), .A2(n5880), .ZN(n1760) );
  OAI21_X1 U1081 ( .B1(n6092), .B2(n1744), .A(n1761), .ZN(n3853) );
  NAND2_X1 U1082 ( .A1(n2814), .A2(n5879), .ZN(n1761) );
  OAI21_X1 U1083 ( .B1(n6093), .B2(n1744), .A(n1762), .ZN(n3852) );
  NAND2_X1 U1084 ( .A1(n2813), .A2(n5880), .ZN(n1762) );
  OAI21_X1 U1085 ( .B1(n5515), .B2(n1744), .A(n1763), .ZN(n3851) );
  NAND2_X1 U1086 ( .A1(n2812), .A2(n5879), .ZN(n1763) );
  OAI21_X1 U1087 ( .B1(n5518), .B2(n1744), .A(n1764), .ZN(n3850) );
  NAND2_X1 U1088 ( .A1(n2811), .A2(n5879), .ZN(n1764) );
  OAI21_X1 U1089 ( .B1(n5521), .B2(n5879), .A(n1765), .ZN(n3849) );
  NAND2_X1 U1090 ( .A1(n2810), .A2(n5880), .ZN(n1765) );
  OAI21_X1 U1091 ( .B1(n5524), .B2(n5880), .A(n1766), .ZN(n3848) );
  NAND2_X1 U1092 ( .A1(n2809), .A2(n5880), .ZN(n1766) );
  OAI21_X1 U1093 ( .B1(n6098), .B2(n5880), .A(n1767), .ZN(n3847) );
  NAND2_X1 U1094 ( .A1(n2808), .A2(n5879), .ZN(n1767) );
  OAI21_X1 U1095 ( .B1(n5530), .B2(n5879), .A(n1768), .ZN(n3846) );
  NAND2_X1 U1096 ( .A1(n2807), .A2(n5880), .ZN(n1768) );
  OAI21_X1 U1097 ( .B1(n5533), .B2(n5880), .A(n1769), .ZN(n3845) );
  NAND2_X1 U1098 ( .A1(n1744), .A2(n6548), .ZN(n1769) );
  OAI21_X1 U1099 ( .B1(n5536), .B2(n5879), .A(n1770), .ZN(n3844) );
  NAND2_X1 U1100 ( .A1(n5880), .A2(n6549), .ZN(n1770) );
  OAI21_X1 U1101 ( .B1(n5539), .B2(n5880), .A(n1771), .ZN(n3843) );
  NAND2_X1 U1102 ( .A1(n5879), .A2(n6550), .ZN(n1771) );
  OAI21_X1 U1103 ( .B1(n5542), .B2(n5879), .A(n1772), .ZN(n3842) );
  NAND2_X1 U1104 ( .A1(n1744), .A2(n6551), .ZN(n1772) );
  OAI21_X1 U1105 ( .B1(n5545), .B2(n5880), .A(n1773), .ZN(n3841) );
  NAND2_X1 U1106 ( .A1(n5880), .A2(n6552), .ZN(n1773) );
  OAI21_X1 U1107 ( .B1(n6105), .B2(n5879), .A(n1774), .ZN(n3840) );
  NAND2_X1 U1108 ( .A1(n5879), .A2(n6553), .ZN(n1774) );
  OAI21_X1 U1109 ( .B1(n5551), .B2(n5880), .A(n1775), .ZN(n3839) );
  NAND2_X1 U1110 ( .A1(n5880), .A2(n6554), .ZN(n1775) );
  OAI21_X1 U1111 ( .B1(n5554), .B2(n1744), .A(n1776), .ZN(n3838) );
  NAND2_X1 U1112 ( .A1(n1744), .A2(n6555), .ZN(n1776) );
  NAND2_X1 U1113 ( .A1(n1777), .A2(n1778), .ZN(n1744) );
  OAI21_X1 U1114 ( .B1(n5461), .B2(n5876), .A(n1780), .ZN(n3837) );
  NAND2_X1 U1115 ( .A1(n1779), .A2(n6556), .ZN(n1780) );
  OAI21_X1 U1116 ( .B1(n6077), .B2(n5876), .A(n1781), .ZN(n3836) );
  NAND2_X1 U1117 ( .A1(n1779), .A2(n6557), .ZN(n1781) );
  OAI21_X1 U1118 ( .B1(n5467), .B2(n5876), .A(n1782), .ZN(n3835) );
  NAND2_X1 U1119 ( .A1(n1779), .A2(n6558), .ZN(n1782) );
  OAI21_X1 U1120 ( .B1(n5470), .B2(n5876), .A(n1783), .ZN(n3834) );
  NAND2_X1 U1121 ( .A1(n1779), .A2(n6559), .ZN(n1783) );
  OAI21_X1 U1122 ( .B1(n5473), .B2(n5876), .A(n1784), .ZN(n3833) );
  NAND2_X1 U1123 ( .A1(n1779), .A2(n6560), .ZN(n1784) );
  OAI21_X1 U1124 ( .B1(n5476), .B2(n5876), .A(n1785), .ZN(n3832) );
  NAND2_X1 U1125 ( .A1(n1779), .A2(n6561), .ZN(n1785) );
  OAI21_X1 U1126 ( .B1(n6082), .B2(n5876), .A(n1786), .ZN(n3831) );
  NAND2_X1 U1127 ( .A1(n1779), .A2(n6562), .ZN(n1786) );
  OAI21_X1 U1128 ( .B1(n5482), .B2(n5876), .A(n1787), .ZN(n3830) );
  NAND2_X1 U1129 ( .A1(n5877), .A2(n6563), .ZN(n1787) );
  OAI21_X1 U1130 ( .B1(n5485), .B2(n5876), .A(n1788), .ZN(n3829) );
  NAND2_X1 U1131 ( .A1(n5876), .A2(n6564), .ZN(n1788) );
  OAI21_X1 U1132 ( .B1(n5488), .B2(n5876), .A(n1789), .ZN(n3828) );
  NAND2_X1 U1133 ( .A1(n5877), .A2(n6565), .ZN(n1789) );
  OAI21_X1 U1134 ( .B1(n5491), .B2(n5876), .A(n1790), .ZN(n3827) );
  NAND2_X1 U1135 ( .A1(n5876), .A2(n6566), .ZN(n1790) );
  OAI21_X1 U1136 ( .B1(n5494), .B2(n5877), .A(n1791), .ZN(n3826) );
  NAND2_X1 U1137 ( .A1(n5877), .A2(n6567), .ZN(n1791) );
  OAI21_X1 U1138 ( .B1(n5497), .B2(n5877), .A(n1792), .ZN(n3825) );
  NAND2_X1 U1139 ( .A1(n5876), .A2(n6568), .ZN(n1792) );
  OAI21_X1 U1140 ( .B1(n5500), .B2(n5877), .A(n1793), .ZN(n3824) );
  NAND2_X1 U1141 ( .A1(n5877), .A2(n6569), .ZN(n1793) );
  OAI21_X1 U1142 ( .B1(n5503), .B2(n5877), .A(n1794), .ZN(n3823) );
  NAND2_X1 U1143 ( .A1(n5876), .A2(n6570), .ZN(n1794) );
  OAI21_X1 U1144 ( .B1(n5506), .B2(n5877), .A(n1795), .ZN(n3822) );
  NAND2_X1 U1145 ( .A1(n1779), .A2(n6571), .ZN(n1795) );
  OAI21_X1 U1146 ( .B1(n6092), .B2(n5877), .A(n1796), .ZN(n3821) );
  NAND2_X1 U1147 ( .A1(n1779), .A2(n6572), .ZN(n1796) );
  OAI21_X1 U1148 ( .B1(n6093), .B2(n5877), .A(n1797), .ZN(n3820) );
  NAND2_X1 U1149 ( .A1(n1779), .A2(n6573), .ZN(n1797) );
  OAI21_X1 U1150 ( .B1(n5515), .B2(n5877), .A(n1798), .ZN(n3819) );
  NAND2_X1 U1151 ( .A1(n1779), .A2(n6574), .ZN(n1798) );
  OAI21_X1 U1152 ( .B1(n5518), .B2(n5877), .A(n1799), .ZN(n3818) );
  NAND2_X1 U1153 ( .A1(n5876), .A2(n6575), .ZN(n1799) );
  OAI21_X1 U1154 ( .B1(n5521), .B2(n5877), .A(n1800), .ZN(n3817) );
  NAND2_X1 U1155 ( .A1(n1779), .A2(n6576), .ZN(n1800) );
  OAI21_X1 U1156 ( .B1(n5524), .B2(n5877), .A(n1801), .ZN(n3816) );
  NAND2_X1 U1157 ( .A1(n1779), .A2(n6577), .ZN(n1801) );
  OAI21_X1 U1158 ( .B1(n6098), .B2(n5877), .A(n1802), .ZN(n3815) );
  NAND2_X1 U1159 ( .A1(n1779), .A2(n6578), .ZN(n1802) );
  OAI21_X1 U1160 ( .B1(n5530), .B2(n5877), .A(n1803), .ZN(n3814) );
  NAND2_X1 U1161 ( .A1(n1779), .A2(n6579), .ZN(n1803) );
  OAI21_X1 U1162 ( .B1(n5533), .B2(n5876), .A(n1804), .ZN(n3813) );
  NAND2_X1 U1163 ( .A1(n1779), .A2(n6580), .ZN(n1804) );
  OAI21_X1 U1164 ( .B1(n5536), .B2(n5877), .A(n1805), .ZN(n3812) );
  NAND2_X1 U1165 ( .A1(n1779), .A2(n6581), .ZN(n1805) );
  OAI21_X1 U1166 ( .B1(n5539), .B2(n5876), .A(n1806), .ZN(n3811) );
  NAND2_X1 U1167 ( .A1(n1779), .A2(n6582), .ZN(n1806) );
  OAI21_X1 U1168 ( .B1(n5542), .B2(n5877), .A(n1807), .ZN(n3810) );
  NAND2_X1 U1169 ( .A1(n1779), .A2(n6583), .ZN(n1807) );
  OAI21_X1 U1170 ( .B1(n5545), .B2(n5876), .A(n1808), .ZN(n3809) );
  NAND2_X1 U1171 ( .A1(n1779), .A2(n6584), .ZN(n1808) );
  OAI21_X1 U1172 ( .B1(n6105), .B2(n5877), .A(n1809), .ZN(n3808) );
  NAND2_X1 U1173 ( .A1(n1779), .A2(n6585), .ZN(n1809) );
  OAI21_X1 U1174 ( .B1(n5551), .B2(n5876), .A(n1810), .ZN(n3807) );
  NAND2_X1 U1175 ( .A1(n1779), .A2(n6586), .ZN(n1810) );
  OAI21_X1 U1176 ( .B1(n5554), .B2(n5877), .A(n1811), .ZN(n3806) );
  NAND2_X1 U1177 ( .A1(n1779), .A2(n6587), .ZN(n1811) );
  NAND2_X1 U1178 ( .A1(n1812), .A2(n1777), .ZN(n1779) );
  OAI21_X1 U1179 ( .B1(n6093), .B2(n5889), .A(n1813), .ZN(n3805) );
  NAND2_X1 U1180 ( .A1(n1726), .A2(n6469), .ZN(n1813) );
  OAI21_X1 U1181 ( .B1(n5515), .B2(n5889), .A(n1814), .ZN(n3804) );
  NAND2_X1 U1182 ( .A1(n1726), .A2(n6470), .ZN(n1814) );
  OAI21_X1 U1183 ( .B1(n5518), .B2(n5889), .A(n1815), .ZN(n3803) );
  NAND2_X1 U1184 ( .A1(n5888), .A2(n6471), .ZN(n1815) );
  OAI21_X1 U1185 ( .B1(n5521), .B2(n5889), .A(n1816), .ZN(n3802) );
  NAND2_X1 U1186 ( .A1(n1726), .A2(n6472), .ZN(n1816) );
  OAI21_X1 U1187 ( .B1(n5524), .B2(n5889), .A(n1817), .ZN(n3801) );
  NAND2_X1 U1188 ( .A1(n1726), .A2(n6473), .ZN(n1817) );
  OAI21_X1 U1189 ( .B1(n6098), .B2(n5889), .A(n1818), .ZN(n3800) );
  NAND2_X1 U1190 ( .A1(n1726), .A2(n6474), .ZN(n1818) );
  OAI21_X1 U1191 ( .B1(n5530), .B2(n5889), .A(n1819), .ZN(n3799) );
  NAND2_X1 U1192 ( .A1(n1726), .A2(n6475), .ZN(n1819) );
  OAI21_X1 U1193 ( .B1(n5533), .B2(n5888), .A(n1820), .ZN(n3798) );
  NAND2_X1 U1194 ( .A1(n1726), .A2(n6476), .ZN(n1820) );
  OAI21_X1 U1195 ( .B1(n5536), .B2(n5889), .A(n1821), .ZN(n3797) );
  NAND2_X1 U1196 ( .A1(n1726), .A2(n6477), .ZN(n1821) );
  OAI21_X1 U1197 ( .B1(n5539), .B2(n5888), .A(n1822), .ZN(n3796) );
  NAND2_X1 U1198 ( .A1(n1726), .A2(n6478), .ZN(n1822) );
  OAI21_X1 U1199 ( .B1(n5542), .B2(n5889), .A(n1823), .ZN(n3795) );
  NAND2_X1 U1200 ( .A1(n1726), .A2(n6479), .ZN(n1823) );
  OAI21_X1 U1201 ( .B1(n5545), .B2(n5888), .A(n1824), .ZN(n3794) );
  NAND2_X1 U1202 ( .A1(n1726), .A2(n6480), .ZN(n1824) );
  OAI21_X1 U1203 ( .B1(n6105), .B2(n5889), .A(n1825), .ZN(n3793) );
  NAND2_X1 U1204 ( .A1(n1726), .A2(n6481), .ZN(n1825) );
  OAI21_X1 U1205 ( .B1(n5551), .B2(n5888), .A(n1826), .ZN(n3792) );
  NAND2_X1 U1206 ( .A1(n1726), .A2(n6482), .ZN(n1826) );
  OAI21_X1 U1207 ( .B1(n5554), .B2(n5889), .A(n1827), .ZN(n3791) );
  NAND2_X1 U1208 ( .A1(n1726), .A2(n6483), .ZN(n1827) );
  NAND2_X1 U1209 ( .A1(n1692), .A2(n1624), .ZN(n1726) );
  OAI21_X1 U1210 ( .B1(n5461), .B2(n5872), .A(n1829), .ZN(n3790) );
  NAND2_X1 U1211 ( .A1(n5872), .A2(n6420), .ZN(n1829) );
  OAI21_X1 U1212 ( .B1(n6077), .B2(n5868), .A(n1830), .ZN(n3789) );
  NAND2_X1 U1213 ( .A1(n1828), .A2(n6421), .ZN(n1830) );
  OAI21_X1 U1214 ( .B1(n5467), .B2(n5872), .A(n1831), .ZN(n3788) );
  NAND2_X1 U1215 ( .A1(n5868), .A2(n6422), .ZN(n1831) );
  OAI21_X1 U1216 ( .B1(n5470), .B2(n5868), .A(n1832), .ZN(n3787) );
  NAND2_X1 U1217 ( .A1(n5872), .A2(n6423), .ZN(n1832) );
  OAI21_X1 U1218 ( .B1(n5473), .B2(n5872), .A(n1833), .ZN(n3786) );
  NAND2_X1 U1219 ( .A1(n5868), .A2(n6424), .ZN(n1833) );
  OAI21_X1 U1220 ( .B1(n5476), .B2(n5868), .A(n1834), .ZN(n3785) );
  NAND2_X1 U1221 ( .A1(n5868), .A2(n6425), .ZN(n1834) );
  OAI21_X1 U1222 ( .B1(n6082), .B2(n5872), .A(n1835), .ZN(n3784) );
  NAND2_X1 U1223 ( .A1(n5868), .A2(n6426), .ZN(n1835) );
  OAI21_X1 U1224 ( .B1(n5482), .B2(n5868), .A(n1836), .ZN(n3783) );
  NAND2_X1 U1225 ( .A1(n1828), .A2(n6427), .ZN(n1836) );
  OAI21_X1 U1226 ( .B1(n5485), .B2(n5872), .A(n1837), .ZN(n3782) );
  NAND2_X1 U1227 ( .A1(n1828), .A2(n6428), .ZN(n1837) );
  OAI21_X1 U1228 ( .B1(n5488), .B2(n5868), .A(n1838), .ZN(n3781) );
  NAND2_X1 U1229 ( .A1(n1828), .A2(n6429), .ZN(n1838) );
  OAI21_X1 U1230 ( .B1(n5491), .B2(n5872), .A(n1839), .ZN(n3780) );
  NAND2_X1 U1231 ( .A1(n1828), .A2(n6430), .ZN(n1839) );
  OAI21_X1 U1232 ( .B1(n5494), .B2(n5872), .A(n1840), .ZN(n3779) );
  NAND2_X1 U1233 ( .A1(n1828), .A2(n6431), .ZN(n1840) );
  OAI21_X1 U1234 ( .B1(n5497), .B2(n5868), .A(n1841), .ZN(n3778) );
  NAND2_X1 U1235 ( .A1(n1828), .A2(n6432), .ZN(n1841) );
  OAI21_X1 U1236 ( .B1(n5500), .B2(n5868), .A(n1842), .ZN(n3777) );
  NAND2_X1 U1237 ( .A1(n1828), .A2(n6433), .ZN(n1842) );
  OAI21_X1 U1238 ( .B1(n5503), .B2(n5872), .A(n1843), .ZN(n3776) );
  NAND2_X1 U1239 ( .A1(n1828), .A2(n6434), .ZN(n1843) );
  OAI21_X1 U1240 ( .B1(n5506), .B2(n5868), .A(n1844), .ZN(n3775) );
  NAND2_X1 U1241 ( .A1(n1828), .A2(n6435), .ZN(n1844) );
  OAI21_X1 U1242 ( .B1(n6092), .B2(n1828), .A(n1845), .ZN(n3774) );
  NAND2_X1 U1243 ( .A1(n5868), .A2(n6436), .ZN(n1845) );
  OAI21_X1 U1244 ( .B1(n5554), .B2(n1846), .A(n1847), .ZN(n3773) );
  NAND2_X1 U1245 ( .A1(n321), .A2(n5861), .ZN(n1847) );
  OAI21_X1 U1246 ( .B1(n5551), .B2(n5863), .A(n1848), .ZN(n3772) );
  NAND2_X1 U1247 ( .A1(n322), .A2(n5861), .ZN(n1848) );
  OAI21_X1 U1248 ( .B1(n6105), .B2(n1846), .A(n1849), .ZN(n3771) );
  NAND2_X1 U1249 ( .A1(n323), .A2(n5861), .ZN(n1849) );
  OAI21_X1 U1250 ( .B1(n5545), .B2(n5861), .A(n1850), .ZN(n3770) );
  NAND2_X1 U1251 ( .A1(n324), .A2(n5861), .ZN(n1850) );
  OAI21_X1 U1252 ( .B1(n5542), .B2(n1846), .A(n1851), .ZN(n3769) );
  NAND2_X1 U1253 ( .A1(n325), .A2(n5861), .ZN(n1851) );
  OAI21_X1 U1254 ( .B1(n5539), .B2(n5863), .A(n1852), .ZN(n3768) );
  NAND2_X1 U1255 ( .A1(n326), .A2(n5863), .ZN(n1852) );
  OAI21_X1 U1256 ( .B1(n5536), .B2(n1846), .A(n1853), .ZN(n3767) );
  NAND2_X1 U1257 ( .A1(n327), .A2(n5863), .ZN(n1853) );
  OAI21_X1 U1258 ( .B1(n5533), .B2(n5861), .A(n1854), .ZN(n3766) );
  NAND2_X1 U1259 ( .A1(n328), .A2(n5863), .ZN(n1854) );
  OAI21_X1 U1260 ( .B1(n5530), .B2(n1846), .A(n1855), .ZN(n3765) );
  NAND2_X1 U1261 ( .A1(n329), .A2(n5863), .ZN(n1855) );
  OAI21_X1 U1262 ( .B1(n6098), .B2(n5861), .A(n1856), .ZN(n3764) );
  NAND2_X1 U1263 ( .A1(n330), .A2(n5863), .ZN(n1856) );
  OAI21_X1 U1264 ( .B1(n5524), .B2(n5863), .A(n1857), .ZN(n3763) );
  NAND2_X1 U1265 ( .A1(n331), .A2(n5863), .ZN(n1857) );
  OAI21_X1 U1266 ( .B1(n5521), .B2(n1846), .A(n1858), .ZN(n3762) );
  NAND2_X1 U1267 ( .A1(n332), .A2(n5863), .ZN(n1858) );
  OAI21_X1 U1268 ( .B1(n5518), .B2(n1846), .A(n1859), .ZN(n3761) );
  NAND2_X1 U1269 ( .A1(n333), .A2(n5863), .ZN(n1859) );
  OAI21_X1 U1270 ( .B1(n5515), .B2(n1846), .A(n1860), .ZN(n3760) );
  NAND2_X1 U1271 ( .A1(n334), .A2(n5863), .ZN(n1860) );
  OAI21_X1 U1272 ( .B1(n6093), .B2(n1846), .A(n1861), .ZN(n3759) );
  NAND2_X1 U1273 ( .A1(n335), .A2(n5863), .ZN(n1861) );
  OAI21_X1 U1274 ( .B1(n6092), .B2(n1846), .A(n1862), .ZN(n3758) );
  NAND2_X1 U1275 ( .A1(n336), .A2(n5863), .ZN(n1862) );
  OAI21_X1 U1276 ( .B1(n6091), .B2(n1846), .A(n1863), .ZN(n3757) );
  NAND2_X1 U1277 ( .A1(n337), .A2(n5861), .ZN(n1863) );
  OAI21_X1 U1278 ( .B1(n5503), .B2(n1846), .A(n1864), .ZN(n3756) );
  NAND2_X1 U1279 ( .A1(n338), .A2(n5863), .ZN(n1864) );
  OAI21_X1 U1280 ( .B1(n6089), .B2(n5861), .A(n1865), .ZN(n3755) );
  NAND2_X1 U1281 ( .A1(n339), .A2(n5861), .ZN(n1865) );
  OAI21_X1 U1282 ( .B1(n6088), .B2(n5863), .A(n1866), .ZN(n3754) );
  NAND2_X1 U1283 ( .A1(n340), .A2(n5863), .ZN(n1866) );
  OAI21_X1 U1284 ( .B1(n6087), .B2(n5863), .A(n1867), .ZN(n3753) );
  NAND2_X1 U1285 ( .A1(n341), .A2(n5863), .ZN(n1867) );
  OAI21_X1 U1286 ( .B1(n6086), .B2(n1846), .A(n1868), .ZN(n3752) );
  NAND2_X1 U1287 ( .A1(n342), .A2(n1846), .ZN(n1868) );
  OAI21_X1 U1288 ( .B1(n6085), .B2(n1846), .A(n1869), .ZN(n3751) );
  NAND2_X1 U1289 ( .A1(n343), .A2(n5861), .ZN(n1869) );
  OAI21_X1 U1290 ( .B1(n6084), .B2(n1846), .A(n1870), .ZN(n3750) );
  NAND2_X1 U1291 ( .A1(n344), .A2(n5863), .ZN(n1870) );
  OAI21_X1 U1292 ( .B1(n6083), .B2(n1846), .A(n1871), .ZN(n3749) );
  NAND2_X1 U1293 ( .A1(n345), .A2(n5861), .ZN(n1871) );
  OAI21_X1 U1294 ( .B1(n6082), .B2(n1846), .A(n1872), .ZN(n3748) );
  NAND2_X1 U1295 ( .A1(n346), .A2(n5861), .ZN(n1872) );
  OAI21_X1 U1296 ( .B1(n6081), .B2(n1846), .A(n1873), .ZN(n3747) );
  NAND2_X1 U1297 ( .A1(n347), .A2(n5861), .ZN(n1873) );
  OAI21_X1 U1298 ( .B1(n6080), .B2(n1846), .A(n1874), .ZN(n3746) );
  NAND2_X1 U1299 ( .A1(n348), .A2(n5861), .ZN(n1874) );
  OAI21_X1 U1300 ( .B1(n6079), .B2(n1846), .A(n1875), .ZN(n3745) );
  NAND2_X1 U1301 ( .A1(n349), .A2(n5861), .ZN(n1875) );
  OAI21_X1 U1302 ( .B1(n6078), .B2(n1846), .A(n1876), .ZN(n3744) );
  NAND2_X1 U1303 ( .A1(n350), .A2(n5861), .ZN(n1876) );
  OAI21_X1 U1304 ( .B1(n5463), .B2(n1846), .A(n1877), .ZN(n3743) );
  NAND2_X1 U1305 ( .A1(n351), .A2(n5861), .ZN(n1877) );
  OAI21_X1 U1306 ( .B1(n6076), .B2(n5863), .A(n1878), .ZN(n3742) );
  NAND2_X1 U1307 ( .A1(n352), .A2(n5861), .ZN(n1878) );
  NAND2_X1 U1308 ( .A1(n1777), .A2(n1658), .ZN(n1846) );
  OAI21_X1 U1309 ( .B1(n5554), .B2(n5860), .A(n1880), .ZN(n3741) );
  NAND2_X1 U1310 ( .A1(n353), .A2(n1879), .ZN(n1880) );
  OAI21_X1 U1311 ( .B1(n6106), .B2(n5859), .A(n1881), .ZN(n3740) );
  NAND2_X1 U1312 ( .A1(n354), .A2(n1879), .ZN(n1881) );
  OAI21_X1 U1313 ( .B1(n5547), .B2(n5860), .A(n1882), .ZN(n3739) );
  NAND2_X1 U1314 ( .A1(n355), .A2(n1879), .ZN(n1882) );
  OAI21_X1 U1315 ( .B1(n6104), .B2(n5859), .A(n1883), .ZN(n3738) );
  NAND2_X1 U1316 ( .A1(n356), .A2(n1879), .ZN(n1883) );
  OAI21_X1 U1317 ( .B1(n6103), .B2(n5860), .A(n1884), .ZN(n3737) );
  NAND2_X1 U1318 ( .A1(n357), .A2(n1879), .ZN(n1884) );
  OAI21_X1 U1319 ( .B1(n6102), .B2(n5859), .A(n1885), .ZN(n3736) );
  NAND2_X1 U1320 ( .A1(n358), .A2(n1879), .ZN(n1885) );
  OAI21_X1 U1321 ( .B1(n6101), .B2(n5860), .A(n1886), .ZN(n3735) );
  NAND2_X1 U1322 ( .A1(n359), .A2(n5860), .ZN(n1886) );
  OAI21_X1 U1323 ( .B1(n6100), .B2(n5859), .A(n1887), .ZN(n3734) );
  NAND2_X1 U1324 ( .A1(n360), .A2(n5859), .ZN(n1887) );
  OAI21_X1 U1325 ( .B1(n6099), .B2(n5860), .A(n1888), .ZN(n3733) );
  NAND2_X1 U1326 ( .A1(n361), .A2(n1879), .ZN(n1888) );
  OAI21_X1 U1327 ( .B1(n6098), .B2(n5859), .A(n1889), .ZN(n3732) );
  NAND2_X1 U1328 ( .A1(n362), .A2(n1879), .ZN(n1889) );
  OAI21_X1 U1329 ( .B1(n6097), .B2(n5860), .A(n1890), .ZN(n3731) );
  NAND2_X1 U1330 ( .A1(n363), .A2(n1879), .ZN(n1890) );
  OAI21_X1 U1331 ( .B1(n6096), .B2(n5859), .A(n1891), .ZN(n3730) );
  NAND2_X1 U1332 ( .A1(n364), .A2(n1879), .ZN(n1891) );
  OAI21_X1 U1333 ( .B1(n6095), .B2(n5859), .A(n1892), .ZN(n3729) );
  NAND2_X1 U1334 ( .A1(n365), .A2(n1879), .ZN(n1892) );
  OAI21_X1 U1335 ( .B1(n6094), .B2(n5859), .A(n1893), .ZN(n3728) );
  NAND2_X1 U1336 ( .A1(n366), .A2(n1879), .ZN(n1893) );
  OAI21_X1 U1337 ( .B1(n5511), .B2(n5859), .A(n1894), .ZN(n3727) );
  NAND2_X1 U1338 ( .A1(n367), .A2(n1879), .ZN(n1894) );
  OAI21_X1 U1339 ( .B1(n6092), .B2(n5859), .A(n1895), .ZN(n3726) );
  NAND2_X1 U1340 ( .A1(n368), .A2(n1879), .ZN(n1895) );
  OAI21_X1 U1341 ( .B1(n6091), .B2(n5859), .A(n1896), .ZN(n3725) );
  NAND2_X1 U1342 ( .A1(n369), .A2(n5860), .ZN(n1896) );
  OAI21_X1 U1343 ( .B1(n5503), .B2(n5859), .A(n1897), .ZN(n3724) );
  NAND2_X1 U1344 ( .A1(n370), .A2(n1879), .ZN(n1897) );
  OAI21_X1 U1345 ( .B1(n6089), .B2(n5859), .A(n1898), .ZN(n3723) );
  NAND2_X1 U1346 ( .A1(n371), .A2(n5859), .ZN(n1898) );
  OAI21_X1 U1347 ( .B1(n6088), .B2(n5859), .A(n1899), .ZN(n3722) );
  NAND2_X1 U1348 ( .A1(n372), .A2(n5859), .ZN(n1899) );
  OAI21_X1 U1349 ( .B1(n6087), .B2(n5859), .A(n1900), .ZN(n3721) );
  NAND2_X1 U1350 ( .A1(n373), .A2(n5860), .ZN(n1900) );
  OAI21_X1 U1351 ( .B1(n6086), .B2(n5859), .A(n1901), .ZN(n3720) );
  NAND2_X1 U1352 ( .A1(n374), .A2(n5860), .ZN(n1901) );
  OAI21_X1 U1353 ( .B1(n6085), .B2(n5860), .A(n1902), .ZN(n3719) );
  NAND2_X1 U1354 ( .A1(n375), .A2(n1879), .ZN(n1902) );
  OAI21_X1 U1355 ( .B1(n6084), .B2(n5860), .A(n1903), .ZN(n3718) );
  NAND2_X1 U1356 ( .A1(n376), .A2(n1879), .ZN(n1903) );
  OAI21_X1 U1357 ( .B1(n6083), .B2(n5860), .A(n1904), .ZN(n3717) );
  NAND2_X1 U1358 ( .A1(n377), .A2(n1879), .ZN(n1904) );
  OAI21_X1 U1359 ( .B1(n6082), .B2(n5860), .A(n1905), .ZN(n3716) );
  NAND2_X1 U1360 ( .A1(n378), .A2(n1879), .ZN(n1905) );
  OAI21_X1 U1361 ( .B1(n6081), .B2(n5860), .A(n1906), .ZN(n3715) );
  NAND2_X1 U1362 ( .A1(n379), .A2(n1879), .ZN(n1906) );
  OAI21_X1 U1363 ( .B1(n6080), .B2(n5860), .A(n1907), .ZN(n3714) );
  NAND2_X1 U1364 ( .A1(n380), .A2(n1879), .ZN(n1907) );
  OAI21_X1 U1365 ( .B1(n6079), .B2(n5860), .A(n1908), .ZN(n3713) );
  NAND2_X1 U1366 ( .A1(n381), .A2(n1879), .ZN(n1908) );
  OAI21_X1 U1367 ( .B1(n6078), .B2(n5860), .A(n1909), .ZN(n3712) );
  NAND2_X1 U1368 ( .A1(n382), .A2(n5860), .ZN(n1909) );
  OAI21_X1 U1369 ( .B1(n5463), .B2(n5860), .A(n1910), .ZN(n3711) );
  NAND2_X1 U1370 ( .A1(n383), .A2(n5859), .ZN(n1910) );
  OAI21_X1 U1371 ( .B1(n6076), .B2(n5860), .A(n1911), .ZN(n3710) );
  NAND2_X1 U1372 ( .A1(n384), .A2(n5859), .ZN(n1911) );
  NAND2_X1 U1373 ( .A1(n1777), .A2(n1624), .ZN(n1879) );
  OAI21_X1 U1374 ( .B1(n5554), .B2(n1912), .A(n1913), .ZN(n3709) );
  NAND2_X1 U1375 ( .A1(n641), .A2(n5849), .ZN(n1913) );
  OAI21_X1 U1376 ( .B1(n6106), .B2(n5851), .A(n1914), .ZN(n3708) );
  NAND2_X1 U1377 ( .A1(n642), .A2(n5849), .ZN(n1914) );
  OAI21_X1 U1378 ( .B1(n5547), .B2(n1912), .A(n1915), .ZN(n3707) );
  NAND2_X1 U1379 ( .A1(n643), .A2(n5849), .ZN(n1915) );
  OAI21_X1 U1380 ( .B1(n6104), .B2(n5849), .A(n1916), .ZN(n3706) );
  NAND2_X1 U1381 ( .A1(n644), .A2(n5849), .ZN(n1916) );
  OAI21_X1 U1382 ( .B1(n6103), .B2(n1912), .A(n1917), .ZN(n3705) );
  NAND2_X1 U1383 ( .A1(n645), .A2(n5849), .ZN(n1917) );
  OAI21_X1 U1384 ( .B1(n6102), .B2(n5851), .A(n1918), .ZN(n3704) );
  NAND2_X1 U1385 ( .A1(n646), .A2(n5851), .ZN(n1918) );
  OAI21_X1 U1386 ( .B1(n6101), .B2(n1912), .A(n1919), .ZN(n3703) );
  NAND2_X1 U1387 ( .A1(n647), .A2(n5851), .ZN(n1919) );
  OAI21_X1 U1388 ( .B1(n6100), .B2(n5849), .A(n1920), .ZN(n3702) );
  NAND2_X1 U1389 ( .A1(n648), .A2(n5851), .ZN(n1920) );
  OAI21_X1 U1390 ( .B1(n6099), .B2(n1912), .A(n1921), .ZN(n3701) );
  NAND2_X1 U1391 ( .A1(n649), .A2(n5851), .ZN(n1921) );
  OAI21_X1 U1392 ( .B1(n6098), .B2(n5849), .A(n1922), .ZN(n3700) );
  NAND2_X1 U1393 ( .A1(n650), .A2(n5851), .ZN(n1922) );
  OAI21_X1 U1394 ( .B1(n6097), .B2(n5851), .A(n1923), .ZN(n3699) );
  NAND2_X1 U1395 ( .A1(n651), .A2(n5851), .ZN(n1923) );
  OAI21_X1 U1396 ( .B1(n6096), .B2(n1912), .A(n1924), .ZN(n3698) );
  NAND2_X1 U1397 ( .A1(n652), .A2(n5851), .ZN(n1924) );
  OAI21_X1 U1398 ( .B1(n6095), .B2(n1912), .A(n1925), .ZN(n3697) );
  NAND2_X1 U1399 ( .A1(n653), .A2(n5851), .ZN(n1925) );
  OAI21_X1 U1400 ( .B1(n6094), .B2(n1912), .A(n1926), .ZN(n3696) );
  NAND2_X1 U1401 ( .A1(n654), .A2(n5851), .ZN(n1926) );
  OAI21_X1 U1402 ( .B1(n5511), .B2(n1912), .A(n1927), .ZN(n3695) );
  NAND2_X1 U1403 ( .A1(n655), .A2(n5851), .ZN(n1927) );
  OAI21_X1 U1404 ( .B1(n6092), .B2(n1912), .A(n1928), .ZN(n3694) );
  NAND2_X1 U1405 ( .A1(n656), .A2(n5851), .ZN(n1928) );
  OAI21_X1 U1406 ( .B1(n5506), .B2(n1912), .A(n1929), .ZN(n3693) );
  NAND2_X1 U1407 ( .A1(n657), .A2(n5849), .ZN(n1929) );
  OAI21_X1 U1408 ( .B1(n5503), .B2(n1912), .A(n1930), .ZN(n3692) );
  NAND2_X1 U1409 ( .A1(n658), .A2(n5851), .ZN(n1930) );
  OAI21_X1 U1410 ( .B1(n5500), .B2(n5849), .A(n1931), .ZN(n3691) );
  NAND2_X1 U1411 ( .A1(n659), .A2(n5849), .ZN(n1931) );
  OAI21_X1 U1412 ( .B1(n5497), .B2(n5851), .A(n1932), .ZN(n3690) );
  NAND2_X1 U1413 ( .A1(n660), .A2(n5851), .ZN(n1932) );
  OAI21_X1 U1414 ( .B1(n5494), .B2(n5851), .A(n1933), .ZN(n3689) );
  NAND2_X1 U1415 ( .A1(n661), .A2(n5851), .ZN(n1933) );
  OAI21_X1 U1416 ( .B1(n5491), .B2(n1912), .A(n1934), .ZN(n3688) );
  NAND2_X1 U1417 ( .A1(n662), .A2(n1912), .ZN(n1934) );
  OAI21_X1 U1418 ( .B1(n5488), .B2(n1912), .A(n1935), .ZN(n3687) );
  NAND2_X1 U1419 ( .A1(n663), .A2(n5849), .ZN(n1935) );
  OAI21_X1 U1420 ( .B1(n5485), .B2(n1912), .A(n1936), .ZN(n3686) );
  NAND2_X1 U1421 ( .A1(n664), .A2(n5851), .ZN(n1936) );
  OAI21_X1 U1422 ( .B1(n5482), .B2(n1912), .A(n1937), .ZN(n3685) );
  NAND2_X1 U1423 ( .A1(n665), .A2(n5849), .ZN(n1937) );
  OAI21_X1 U1424 ( .B1(n6082), .B2(n1912), .A(n1938), .ZN(n3684) );
  NAND2_X1 U1425 ( .A1(n666), .A2(n5849), .ZN(n1938) );
  OAI21_X1 U1426 ( .B1(n5476), .B2(n1912), .A(n1939), .ZN(n3683) );
  NAND2_X1 U1427 ( .A1(n667), .A2(n5849), .ZN(n1939) );
  OAI21_X1 U1428 ( .B1(n5473), .B2(n1912), .A(n1940), .ZN(n3682) );
  NAND2_X1 U1429 ( .A1(n668), .A2(n5849), .ZN(n1940) );
  OAI21_X1 U1430 ( .B1(n5470), .B2(n1912), .A(n1941), .ZN(n3681) );
  NAND2_X1 U1431 ( .A1(n669), .A2(n5849), .ZN(n1941) );
  OAI21_X1 U1432 ( .B1(n5467), .B2(n1912), .A(n1942), .ZN(n3680) );
  NAND2_X1 U1433 ( .A1(n670), .A2(n5849), .ZN(n1942) );
  OAI21_X1 U1434 ( .B1(n5463), .B2(n1912), .A(n1943), .ZN(n3679) );
  NAND2_X1 U1435 ( .A1(n671), .A2(n5849), .ZN(n1943) );
  OAI21_X1 U1436 ( .B1(n5461), .B2(n5851), .A(n1944), .ZN(n3678) );
  NAND2_X1 U1437 ( .A1(n672), .A2(n5849), .ZN(n1944) );
  NAND2_X1 U1438 ( .A1(n1777), .A2(n1590), .ZN(n1912) );
  OAI21_X1 U1439 ( .B1(n5554), .B2(n5846), .A(n1946), .ZN(n3677) );
  NAND2_X1 U1440 ( .A1(n481), .A2(n1945), .ZN(n1946) );
  OAI21_X1 U1441 ( .B1(n5551), .B2(n5846), .A(n1947), .ZN(n3676) );
  NAND2_X1 U1442 ( .A1(n482), .A2(n1945), .ZN(n1947) );
  OAI21_X1 U1443 ( .B1(n5547), .B2(n5846), .A(n1948), .ZN(n3675) );
  NAND2_X1 U1444 ( .A1(n483), .A2(n1945), .ZN(n1948) );
  OAI21_X1 U1445 ( .B1(n5545), .B2(n5846), .A(n1949), .ZN(n3674) );
  NAND2_X1 U1446 ( .A1(n484), .A2(n1945), .ZN(n1949) );
  OAI21_X1 U1447 ( .B1(n5542), .B2(n5846), .A(n1950), .ZN(n3673) );
  NAND2_X1 U1448 ( .A1(n485), .A2(n1945), .ZN(n1950) );
  OAI21_X1 U1449 ( .B1(n5539), .B2(n5846), .A(n1951), .ZN(n3672) );
  NAND2_X1 U1450 ( .A1(n486), .A2(n1945), .ZN(n1951) );
  OAI21_X1 U1451 ( .B1(n5536), .B2(n5846), .A(n1952), .ZN(n3671) );
  NAND2_X1 U1452 ( .A1(n487), .A2(n1945), .ZN(n1952) );
  OAI21_X1 U1453 ( .B1(n5533), .B2(n5846), .A(n1953), .ZN(n3670) );
  NAND2_X1 U1454 ( .A1(n488), .A2(n5847), .ZN(n1953) );
  OAI21_X1 U1455 ( .B1(n5530), .B2(n5846), .A(n1954), .ZN(n3669) );
  NAND2_X1 U1456 ( .A1(n489), .A2(n5846), .ZN(n1954) );
  OAI21_X1 U1457 ( .B1(n6098), .B2(n5846), .A(n1955), .ZN(n3668) );
  NAND2_X1 U1458 ( .A1(n490), .A2(n1945), .ZN(n1955) );
  OAI21_X1 U1459 ( .B1(n5524), .B2(n5846), .A(n1956), .ZN(n3667) );
  NAND2_X1 U1460 ( .A1(n491), .A2(n1945), .ZN(n1956) );
  OAI21_X1 U1461 ( .B1(n5521), .B2(n5847), .A(n1957), .ZN(n3666) );
  NAND2_X1 U1462 ( .A1(n492), .A2(n5847), .ZN(n1957) );
  OAI21_X1 U1463 ( .B1(n5518), .B2(n5847), .A(n1958), .ZN(n3665) );
  NAND2_X1 U1464 ( .A1(n493), .A2(n5846), .ZN(n1958) );
  OAI21_X1 U1465 ( .B1(n5515), .B2(n5847), .A(n1959), .ZN(n3664) );
  NAND2_X1 U1466 ( .A1(n494), .A2(n5847), .ZN(n1959) );
  OAI21_X1 U1467 ( .B1(n5511), .B2(n5847), .A(n1960), .ZN(n3663) );
  NAND2_X1 U1468 ( .A1(n495), .A2(n5846), .ZN(n1960) );
  OAI21_X1 U1469 ( .B1(n6092), .B2(n5847), .A(n1961), .ZN(n3662) );
  NAND2_X1 U1470 ( .A1(n496), .A2(n5847), .ZN(n1961) );
  OAI21_X1 U1471 ( .B1(n5506), .B2(n5847), .A(n1962), .ZN(n3661) );
  NAND2_X1 U1472 ( .A1(n497), .A2(n1945), .ZN(n1962) );
  OAI21_X1 U1473 ( .B1(n5503), .B2(n5847), .A(n1963), .ZN(n3660) );
  NAND2_X1 U1474 ( .A1(n498), .A2(n5846), .ZN(n1963) );
  OAI21_X1 U1475 ( .B1(n5500), .B2(n5847), .A(n1964), .ZN(n3659) );
  NAND2_X1 U1476 ( .A1(n499), .A2(n1945), .ZN(n1964) );
  OAI21_X1 U1477 ( .B1(n5497), .B2(n5847), .A(n1965), .ZN(n3658) );
  NAND2_X1 U1478 ( .A1(n500), .A2(n5847), .ZN(n1965) );
  OAI21_X1 U1479 ( .B1(n5494), .B2(n5847), .A(n1966), .ZN(n3657) );
  NAND2_X1 U1480 ( .A1(n501), .A2(n1945), .ZN(n1966) );
  OAI21_X1 U1481 ( .B1(n5491), .B2(n5847), .A(n1967), .ZN(n3656) );
  NAND2_X1 U1482 ( .A1(n502), .A2(n5846), .ZN(n1967) );
  OAI21_X1 U1483 ( .B1(n5488), .B2(n5847), .A(n1968), .ZN(n3655) );
  NAND2_X1 U1484 ( .A1(n503), .A2(n1945), .ZN(n1968) );
  OAI21_X1 U1485 ( .B1(n5485), .B2(n5846), .A(n1969), .ZN(n3654) );
  NAND2_X1 U1486 ( .A1(n504), .A2(n1945), .ZN(n1969) );
  OAI21_X1 U1487 ( .B1(n5482), .B2(n5847), .A(n1970), .ZN(n3653) );
  NAND2_X1 U1488 ( .A1(n505), .A2(n1945), .ZN(n1970) );
  OAI21_X1 U1489 ( .B1(n6082), .B2(n5846), .A(n1971), .ZN(n3652) );
  NAND2_X1 U1490 ( .A1(n506), .A2(n1945), .ZN(n1971) );
  OAI21_X1 U1491 ( .B1(n5476), .B2(n5847), .A(n1972), .ZN(n3651) );
  NAND2_X1 U1492 ( .A1(n507), .A2(n1945), .ZN(n1972) );
  OAI21_X1 U1493 ( .B1(n5473), .B2(n5846), .A(n1973), .ZN(n3650) );
  NAND2_X1 U1494 ( .A1(n508), .A2(n1945), .ZN(n1973) );
  OAI21_X1 U1495 ( .B1(n5470), .B2(n5847), .A(n1974), .ZN(n3649) );
  NAND2_X1 U1496 ( .A1(n509), .A2(n1945), .ZN(n1974) );
  OAI21_X1 U1497 ( .B1(n5467), .B2(n5846), .A(n1975), .ZN(n3648) );
  NAND2_X1 U1498 ( .A1(n510), .A2(n1945), .ZN(n1975) );
  OAI21_X1 U1499 ( .B1(n5463), .B2(n5847), .A(n1976), .ZN(n3647) );
  NAND2_X1 U1500 ( .A1(n511), .A2(n1945), .ZN(n1976) );
  OAI21_X1 U1501 ( .B1(n5461), .B2(n5846), .A(n1977), .ZN(n3646) );
  NAND2_X1 U1502 ( .A1(n512), .A2(n1945), .ZN(n1977) );
  NAND2_X1 U1503 ( .A1(n1777), .A2(n1555), .ZN(n1945) );
  OAI21_X1 U1504 ( .B1(n5554), .B2(n5840), .A(n1979), .ZN(n3645) );
  NAND2_X1 U1505 ( .A1(n513), .A2(n1978), .ZN(n1979) );
  OAI21_X1 U1506 ( .B1(n5551), .B2(n5840), .A(n1980), .ZN(n3644) );
  NAND2_X1 U1507 ( .A1(n514), .A2(n1978), .ZN(n1980) );
  OAI21_X1 U1508 ( .B1(n5547), .B2(n5840), .A(n1981), .ZN(n3643) );
  NAND2_X1 U1509 ( .A1(n515), .A2(n1978), .ZN(n1981) );
  OAI21_X1 U1510 ( .B1(n5545), .B2(n5840), .A(n1982), .ZN(n3642) );
  NAND2_X1 U1511 ( .A1(n516), .A2(n1978), .ZN(n1982) );
  OAI21_X1 U1512 ( .B1(n5542), .B2(n5840), .A(n1983), .ZN(n3641) );
  NAND2_X1 U1513 ( .A1(n517), .A2(n1978), .ZN(n1983) );
  OAI21_X1 U1514 ( .B1(n5539), .B2(n5840), .A(n1984), .ZN(n3640) );
  NAND2_X1 U1515 ( .A1(n518), .A2(n1978), .ZN(n1984) );
  OAI21_X1 U1516 ( .B1(n5536), .B2(n5840), .A(n1985), .ZN(n3639) );
  NAND2_X1 U1517 ( .A1(n519), .A2(n1978), .ZN(n1985) );
  OAI21_X1 U1518 ( .B1(n5533), .B2(n5840), .A(n1986), .ZN(n3638) );
  NAND2_X1 U1519 ( .A1(n520), .A2(n5841), .ZN(n1986) );
  OAI21_X1 U1520 ( .B1(n5530), .B2(n5840), .A(n1987), .ZN(n3637) );
  NAND2_X1 U1521 ( .A1(n521), .A2(n5840), .ZN(n1987) );
  OAI21_X1 U1522 ( .B1(n6098), .B2(n5840), .A(n1988), .ZN(n3636) );
  NAND2_X1 U1523 ( .A1(n522), .A2(n1978), .ZN(n1988) );
  OAI21_X1 U1524 ( .B1(n5524), .B2(n5840), .A(n1989), .ZN(n3635) );
  NAND2_X1 U1525 ( .A1(n523), .A2(n1978), .ZN(n1989) );
  OAI21_X1 U1526 ( .B1(n5521), .B2(n5841), .A(n1990), .ZN(n3634) );
  NAND2_X1 U1527 ( .A1(n524), .A2(n5841), .ZN(n1990) );
  OAI21_X1 U1528 ( .B1(n5518), .B2(n5841), .A(n1991), .ZN(n3633) );
  NAND2_X1 U1529 ( .A1(n525), .A2(n5840), .ZN(n1991) );
  OAI21_X1 U1530 ( .B1(n5515), .B2(n5841), .A(n1992), .ZN(n3632) );
  NAND2_X1 U1531 ( .A1(n526), .A2(n5841), .ZN(n1992) );
  OAI21_X1 U1532 ( .B1(n5511), .B2(n5841), .A(n1993), .ZN(n3631) );
  NAND2_X1 U1533 ( .A1(n527), .A2(n5840), .ZN(n1993) );
  OAI21_X1 U1534 ( .B1(n6092), .B2(n5841), .A(n1994), .ZN(n3630) );
  NAND2_X1 U1535 ( .A1(n528), .A2(n5841), .ZN(n1994) );
  OAI21_X1 U1536 ( .B1(n5506), .B2(n5841), .A(n1995), .ZN(n3629) );
  NAND2_X1 U1537 ( .A1(n529), .A2(n1978), .ZN(n1995) );
  OAI21_X1 U1538 ( .B1(n5503), .B2(n5841), .A(n1996), .ZN(n3628) );
  NAND2_X1 U1539 ( .A1(n530), .A2(n5840), .ZN(n1996) );
  OAI21_X1 U1540 ( .B1(n5500), .B2(n5841), .A(n1997), .ZN(n3627) );
  NAND2_X1 U1541 ( .A1(n531), .A2(n1978), .ZN(n1997) );
  OAI21_X1 U1542 ( .B1(n5497), .B2(n5841), .A(n1998), .ZN(n3626) );
  NAND2_X1 U1543 ( .A1(n532), .A2(n5841), .ZN(n1998) );
  OAI21_X1 U1544 ( .B1(n5494), .B2(n5841), .A(n1999), .ZN(n3625) );
  NAND2_X1 U1545 ( .A1(n533), .A2(n1978), .ZN(n1999) );
  OAI21_X1 U1546 ( .B1(n5491), .B2(n5841), .A(n2000), .ZN(n3624) );
  NAND2_X1 U1547 ( .A1(n534), .A2(n5840), .ZN(n2000) );
  OAI21_X1 U1548 ( .B1(n5488), .B2(n5841), .A(n2001), .ZN(n3623) );
  NAND2_X1 U1549 ( .A1(n535), .A2(n1978), .ZN(n2001) );
  OAI21_X1 U1550 ( .B1(n5485), .B2(n5840), .A(n2002), .ZN(n3622) );
  NAND2_X1 U1551 ( .A1(n536), .A2(n1978), .ZN(n2002) );
  OAI21_X1 U1552 ( .B1(n5482), .B2(n5841), .A(n2003), .ZN(n3621) );
  NAND2_X1 U1553 ( .A1(n537), .A2(n1978), .ZN(n2003) );
  OAI21_X1 U1554 ( .B1(n6082), .B2(n5840), .A(n2004), .ZN(n3620) );
  NAND2_X1 U1555 ( .A1(n538), .A2(n1978), .ZN(n2004) );
  OAI21_X1 U1556 ( .B1(n5476), .B2(n5841), .A(n2005), .ZN(n3619) );
  NAND2_X1 U1557 ( .A1(n539), .A2(n1978), .ZN(n2005) );
  OAI21_X1 U1558 ( .B1(n5473), .B2(n5840), .A(n2006), .ZN(n3618) );
  NAND2_X1 U1559 ( .A1(n540), .A2(n1978), .ZN(n2006) );
  OAI21_X1 U1560 ( .B1(n5470), .B2(n5841), .A(n2007), .ZN(n3617) );
  NAND2_X1 U1561 ( .A1(n541), .A2(n1978), .ZN(n2007) );
  OAI21_X1 U1562 ( .B1(n5467), .B2(n5840), .A(n2008), .ZN(n3616) );
  NAND2_X1 U1563 ( .A1(n542), .A2(n1978), .ZN(n2008) );
  OAI21_X1 U1564 ( .B1(n5463), .B2(n5841), .A(n2009), .ZN(n3615) );
  NAND2_X1 U1565 ( .A1(n543), .A2(n1978), .ZN(n2009) );
  OAI21_X1 U1566 ( .B1(n5461), .B2(n5840), .A(n2010), .ZN(n3614) );
  NAND2_X1 U1567 ( .A1(n544), .A2(n1978), .ZN(n2010) );
  NAND2_X1 U1568 ( .A1(n1692), .A2(n1521), .ZN(n1978) );
  OAI21_X1 U1569 ( .B1(n5554), .B2(n5836), .A(n2012), .ZN(n3613) );
  NAND2_X1 U1570 ( .A1(n705), .A2(n2011), .ZN(n2012) );
  OAI21_X1 U1571 ( .B1(n5551), .B2(n5835), .A(n2013), .ZN(n3612) );
  NAND2_X1 U1572 ( .A1(n706), .A2(n2011), .ZN(n2013) );
  OAI21_X1 U1573 ( .B1(n5547), .B2(n5836), .A(n2014), .ZN(n3611) );
  NAND2_X1 U1574 ( .A1(n707), .A2(n2011), .ZN(n2014) );
  OAI21_X1 U1575 ( .B1(n5545), .B2(n5835), .A(n2015), .ZN(n3610) );
  NAND2_X1 U1576 ( .A1(n708), .A2(n2011), .ZN(n2015) );
  OAI21_X1 U1577 ( .B1(n5542), .B2(n5836), .A(n2016), .ZN(n3609) );
  NAND2_X1 U1578 ( .A1(n709), .A2(n2011), .ZN(n2016) );
  OAI21_X1 U1579 ( .B1(n5539), .B2(n5835), .A(n2017), .ZN(n3608) );
  NAND2_X1 U1580 ( .A1(n710), .A2(n2011), .ZN(n2017) );
  OAI21_X1 U1581 ( .B1(n5536), .B2(n5836), .A(n2018), .ZN(n3607) );
  NAND2_X1 U1582 ( .A1(n711), .A2(n5836), .ZN(n2018) );
  OAI21_X1 U1583 ( .B1(n5533), .B2(n5835), .A(n2019), .ZN(n3606) );
  NAND2_X1 U1584 ( .A1(n712), .A2(n5835), .ZN(n2019) );
  OAI21_X1 U1585 ( .B1(n5530), .B2(n5836), .A(n2020), .ZN(n3605) );
  NAND2_X1 U1586 ( .A1(n713), .A2(n2011), .ZN(n2020) );
  OAI21_X1 U1587 ( .B1(n6098), .B2(n5835), .A(n2021), .ZN(n3604) );
  NAND2_X1 U1588 ( .A1(n714), .A2(n2011), .ZN(n2021) );
  OAI21_X1 U1589 ( .B1(n5524), .B2(n5836), .A(n2022), .ZN(n3603) );
  NAND2_X1 U1590 ( .A1(n715), .A2(n2011), .ZN(n2022) );
  OAI21_X1 U1591 ( .B1(n5521), .B2(n5835), .A(n2023), .ZN(n3602) );
  NAND2_X1 U1592 ( .A1(n716), .A2(n2011), .ZN(n2023) );
  OAI21_X1 U1593 ( .B1(n5518), .B2(n5835), .A(n2024), .ZN(n3601) );
  NAND2_X1 U1594 ( .A1(n717), .A2(n2011), .ZN(n2024) );
  OAI21_X1 U1595 ( .B1(n5515), .B2(n5835), .A(n2025), .ZN(n3600) );
  NAND2_X1 U1596 ( .A1(n718), .A2(n2011), .ZN(n2025) );
  OAI21_X1 U1597 ( .B1(n5511), .B2(n5835), .A(n2026), .ZN(n3599) );
  NAND2_X1 U1598 ( .A1(n719), .A2(n2011), .ZN(n2026) );
  OAI21_X1 U1599 ( .B1(n6092), .B2(n5835), .A(n2027), .ZN(n3598) );
  NAND2_X1 U1600 ( .A1(n720), .A2(n2011), .ZN(n2027) );
  OAI21_X1 U1601 ( .B1(n5506), .B2(n5835), .A(n2028), .ZN(n3597) );
  NAND2_X1 U1602 ( .A1(n721), .A2(n5836), .ZN(n2028) );
  OAI21_X1 U1603 ( .B1(n5503), .B2(n5835), .A(n2029), .ZN(n3596) );
  NAND2_X1 U1604 ( .A1(n722), .A2(n2011), .ZN(n2029) );
  OAI21_X1 U1605 ( .B1(n5500), .B2(n5835), .A(n2030), .ZN(n3595) );
  NAND2_X1 U1606 ( .A1(n723), .A2(n5835), .ZN(n2030) );
  OAI21_X1 U1607 ( .B1(n5497), .B2(n5835), .A(n2031), .ZN(n3594) );
  NAND2_X1 U1608 ( .A1(n724), .A2(n5835), .ZN(n2031) );
  OAI21_X1 U1609 ( .B1(n5494), .B2(n5835), .A(n2032), .ZN(n3593) );
  NAND2_X1 U1610 ( .A1(n725), .A2(n5836), .ZN(n2032) );
  OAI21_X1 U1611 ( .B1(n5491), .B2(n5835), .A(n2033), .ZN(n3592) );
  NAND2_X1 U1612 ( .A1(n726), .A2(n5836), .ZN(n2033) );
  OAI21_X1 U1613 ( .B1(n5488), .B2(n5836), .A(n2034), .ZN(n3591) );
  NAND2_X1 U1614 ( .A1(n727), .A2(n2011), .ZN(n2034) );
  OAI21_X1 U1615 ( .B1(n5485), .B2(n5836), .A(n2035), .ZN(n3590) );
  NAND2_X1 U1616 ( .A1(n728), .A2(n2011), .ZN(n2035) );
  OAI21_X1 U1617 ( .B1(n5482), .B2(n5836), .A(n2036), .ZN(n3589) );
  NAND2_X1 U1618 ( .A1(n729), .A2(n2011), .ZN(n2036) );
  OAI21_X1 U1619 ( .B1(n6082), .B2(n5836), .A(n2037), .ZN(n3588) );
  NAND2_X1 U1620 ( .A1(n730), .A2(n2011), .ZN(n2037) );
  OAI21_X1 U1621 ( .B1(n5476), .B2(n5836), .A(n2038), .ZN(n3587) );
  NAND2_X1 U1622 ( .A1(n731), .A2(n2011), .ZN(n2038) );
  OAI21_X1 U1623 ( .B1(n5473), .B2(n5836), .A(n2039), .ZN(n3586) );
  NAND2_X1 U1624 ( .A1(n732), .A2(n2011), .ZN(n2039) );
  OAI21_X1 U1625 ( .B1(n5470), .B2(n5836), .A(n2040), .ZN(n3585) );
  NAND2_X1 U1626 ( .A1(n733), .A2(n2011), .ZN(n2040) );
  OAI21_X1 U1627 ( .B1(n5467), .B2(n5836), .A(n2041), .ZN(n3584) );
  NAND2_X1 U1628 ( .A1(n734), .A2(n5836), .ZN(n2041) );
  OAI21_X1 U1629 ( .B1(n5463), .B2(n5836), .A(n2042), .ZN(n3583) );
  NAND2_X1 U1630 ( .A1(n735), .A2(n5835), .ZN(n2042) );
  OAI21_X1 U1631 ( .B1(n5461), .B2(n5836), .A(n2043), .ZN(n3582) );
  NAND2_X1 U1632 ( .A1(n736), .A2(n5835), .ZN(n2043) );
  NAND2_X1 U1633 ( .A1(n1812), .A2(n1692), .ZN(n2011) );
  OAI21_X1 U1634 ( .B1(n5554), .B2(n5829), .A(n2045), .ZN(n3581) );
  NAND2_X1 U1635 ( .A1(n2044), .A2(n6387), .ZN(n2045) );
  OAI21_X1 U1636 ( .B1(n5551), .B2(n5830), .A(n2046), .ZN(n3580) );
  NAND2_X1 U1637 ( .A1(n2044), .A2(n6386), .ZN(n2046) );
  OAI21_X1 U1638 ( .B1(n5547), .B2(n5829), .A(n2047), .ZN(n3579) );
  NAND2_X1 U1639 ( .A1(n2044), .A2(n6385), .ZN(n2047) );
  OAI21_X1 U1640 ( .B1(n5545), .B2(n5830), .A(n2048), .ZN(n3578) );
  NAND2_X1 U1641 ( .A1(n2044), .A2(n6384), .ZN(n2048) );
  OAI21_X1 U1642 ( .B1(n5542), .B2(n5829), .A(n2049), .ZN(n3577) );
  NAND2_X1 U1643 ( .A1(n2044), .A2(n6383), .ZN(n2049) );
  OAI21_X1 U1644 ( .B1(n5539), .B2(n5830), .A(n2050), .ZN(n3576) );
  NAND2_X1 U1645 ( .A1(n2044), .A2(n6382), .ZN(n2050) );
  OAI21_X1 U1646 ( .B1(n5536), .B2(n5829), .A(n2051), .ZN(n3575) );
  NAND2_X1 U1647 ( .A1(n5829), .A2(n6381), .ZN(n2051) );
  OAI21_X1 U1648 ( .B1(n5533), .B2(n5830), .A(n2052), .ZN(n3574) );
  NAND2_X1 U1649 ( .A1(n5829), .A2(n6380), .ZN(n2052) );
  OAI21_X1 U1650 ( .B1(n5530), .B2(n5829), .A(n2053), .ZN(n3573) );
  NAND2_X1 U1651 ( .A1(n5830), .A2(n6379), .ZN(n2053) );
  OAI21_X1 U1652 ( .B1(n6098), .B2(n5830), .A(n2054), .ZN(n3572) );
  NAND2_X1 U1653 ( .A1(n2044), .A2(n6378), .ZN(n2054) );
  OAI21_X1 U1654 ( .B1(n5524), .B2(n5829), .A(n2055), .ZN(n3571) );
  NAND2_X1 U1655 ( .A1(n5829), .A2(n6377), .ZN(n2055) );
  OAI21_X1 U1656 ( .B1(n5521), .B2(n5829), .A(n2056), .ZN(n3570) );
  NAND2_X1 U1657 ( .A1(n2044), .A2(n6376), .ZN(n2056) );
  OAI21_X1 U1658 ( .B1(n5518), .B2(n5829), .A(n2057), .ZN(n3569) );
  NAND2_X1 U1659 ( .A1(n2044), .A2(n6375), .ZN(n2057) );
  OAI21_X1 U1660 ( .B1(n5515), .B2(n5829), .A(n2058), .ZN(n3568) );
  NAND2_X1 U1661 ( .A1(n2044), .A2(n6374), .ZN(n2058) );
  OAI21_X1 U1662 ( .B1(n5511), .B2(n5829), .A(n2059), .ZN(n3567) );
  NAND2_X1 U1663 ( .A1(n2044), .A2(n6373), .ZN(n2059) );
  OAI21_X1 U1664 ( .B1(n6092), .B2(n5829), .A(n2060), .ZN(n3566) );
  NAND2_X1 U1665 ( .A1(n2044), .A2(n6372), .ZN(n2060) );
  OAI21_X1 U1666 ( .B1(n5506), .B2(n5829), .A(n2061), .ZN(n3565) );
  NAND2_X1 U1667 ( .A1(n5830), .A2(n6371), .ZN(n2061) );
  OAI21_X1 U1668 ( .B1(n5503), .B2(n5829), .A(n2062), .ZN(n3564) );
  NAND2_X1 U1669 ( .A1(n2044), .A2(n6370), .ZN(n2062) );
  OAI21_X1 U1670 ( .B1(n5500), .B2(n5829), .A(n2063), .ZN(n3563) );
  NAND2_X1 U1671 ( .A1(n5830), .A2(n6369), .ZN(n2063) );
  OAI21_X1 U1672 ( .B1(n5497), .B2(n5829), .A(n2064), .ZN(n3562) );
  NAND2_X1 U1673 ( .A1(n5829), .A2(n6368), .ZN(n2064) );
  OAI21_X1 U1674 ( .B1(n5494), .B2(n5829), .A(n2065), .ZN(n3561) );
  NAND2_X1 U1675 ( .A1(n5830), .A2(n6367), .ZN(n2065) );
  OAI21_X1 U1676 ( .B1(n5491), .B2(n5829), .A(n2066), .ZN(n3560) );
  NAND2_X1 U1677 ( .A1(n5830), .A2(n6366), .ZN(n2066) );
  OAI21_X1 U1678 ( .B1(n5488), .B2(n5830), .A(n2067), .ZN(n3559) );
  NAND2_X1 U1679 ( .A1(n2044), .A2(n6365), .ZN(n2067) );
  OAI21_X1 U1680 ( .B1(n5485), .B2(n5830), .A(n2068), .ZN(n3558) );
  NAND2_X1 U1681 ( .A1(n2044), .A2(n6364), .ZN(n2068) );
  OAI21_X1 U1682 ( .B1(n5482), .B2(n5830), .A(n2069), .ZN(n3557) );
  NAND2_X1 U1683 ( .A1(n2044), .A2(n6363), .ZN(n2069) );
  OAI21_X1 U1684 ( .B1(n6082), .B2(n5830), .A(n2070), .ZN(n3556) );
  NAND2_X1 U1685 ( .A1(n2044), .A2(n6362), .ZN(n2070) );
  OAI21_X1 U1686 ( .B1(n5476), .B2(n5830), .A(n2071), .ZN(n3555) );
  NAND2_X1 U1687 ( .A1(n2044), .A2(n6361), .ZN(n2071) );
  OAI21_X1 U1688 ( .B1(n5473), .B2(n5830), .A(n2072), .ZN(n3554) );
  NAND2_X1 U1689 ( .A1(n2044), .A2(n6360), .ZN(n2072) );
  OAI21_X1 U1690 ( .B1(n5470), .B2(n5830), .A(n2073), .ZN(n3553) );
  NAND2_X1 U1691 ( .A1(n2044), .A2(n6359), .ZN(n2073) );
  OAI21_X1 U1692 ( .B1(n5467), .B2(n5830), .A(n2074), .ZN(n3552) );
  NAND2_X1 U1693 ( .A1(n2044), .A2(n6358), .ZN(n2074) );
  OAI21_X1 U1694 ( .B1(n5463), .B2(n5830), .A(n2075), .ZN(n3551) );
  NAND2_X1 U1695 ( .A1(n2044), .A2(n6357), .ZN(n2075) );
  OAI21_X1 U1696 ( .B1(n5461), .B2(n5830), .A(n2076), .ZN(n3550) );
  NAND2_X1 U1697 ( .A1(n2044), .A2(n6356), .ZN(n2076) );
  NAND2_X1 U1698 ( .A1(n1778), .A2(n1692), .ZN(n2044) );
  OAI21_X1 U1699 ( .B1(n5554), .B2(n2077), .A(n2078), .ZN(n3549) );
  NAND2_X1 U1700 ( .A1(n673), .A2(n5819), .ZN(n2078) );
  OAI21_X1 U1701 ( .B1(n5551), .B2(n5821), .A(n2079), .ZN(n3548) );
  NAND2_X1 U1702 ( .A1(n674), .A2(n5819), .ZN(n2079) );
  OAI21_X1 U1703 ( .B1(n5547), .B2(n2077), .A(n2080), .ZN(n3547) );
  NAND2_X1 U1704 ( .A1(n675), .A2(n5819), .ZN(n2080) );
  OAI21_X1 U1705 ( .B1(n5545), .B2(n5819), .A(n2081), .ZN(n3546) );
  NAND2_X1 U1706 ( .A1(n676), .A2(n5819), .ZN(n2081) );
  OAI21_X1 U1707 ( .B1(n5542), .B2(n2077), .A(n2082), .ZN(n3545) );
  NAND2_X1 U1708 ( .A1(n677), .A2(n5819), .ZN(n2082) );
  OAI21_X1 U1709 ( .B1(n5539), .B2(n5821), .A(n2083), .ZN(n3544) );
  NAND2_X1 U1710 ( .A1(n678), .A2(n5821), .ZN(n2083) );
  OAI21_X1 U1711 ( .B1(n5536), .B2(n2077), .A(n2084), .ZN(n3543) );
  NAND2_X1 U1712 ( .A1(n679), .A2(n5821), .ZN(n2084) );
  OAI21_X1 U1713 ( .B1(n5533), .B2(n5819), .A(n2085), .ZN(n3542) );
  NAND2_X1 U1714 ( .A1(n680), .A2(n5821), .ZN(n2085) );
  OAI21_X1 U1715 ( .B1(n5530), .B2(n2077), .A(n2086), .ZN(n3541) );
  NAND2_X1 U1716 ( .A1(n681), .A2(n5821), .ZN(n2086) );
  OAI21_X1 U1717 ( .B1(n6098), .B2(n5819), .A(n2087), .ZN(n3540) );
  NAND2_X1 U1718 ( .A1(n682), .A2(n5821), .ZN(n2087) );
  OAI21_X1 U1719 ( .B1(n5524), .B2(n5821), .A(n2088), .ZN(n3539) );
  NAND2_X1 U1720 ( .A1(n683), .A2(n5821), .ZN(n2088) );
  OAI21_X1 U1721 ( .B1(n5521), .B2(n2077), .A(n2089), .ZN(n3538) );
  NAND2_X1 U1722 ( .A1(n684), .A2(n5821), .ZN(n2089) );
  OAI21_X1 U1723 ( .B1(n5518), .B2(n2077), .A(n2090), .ZN(n3537) );
  NAND2_X1 U1724 ( .A1(n685), .A2(n5821), .ZN(n2090) );
  OAI21_X1 U1725 ( .B1(n5515), .B2(n2077), .A(n2091), .ZN(n3536) );
  NAND2_X1 U1726 ( .A1(n686), .A2(n5821), .ZN(n2091) );
  OAI21_X1 U1727 ( .B1(n5511), .B2(n2077), .A(n2092), .ZN(n3535) );
  NAND2_X1 U1728 ( .A1(n687), .A2(n5821), .ZN(n2092) );
  OAI21_X1 U1729 ( .B1(n6092), .B2(n2077), .A(n2093), .ZN(n3534) );
  NAND2_X1 U1730 ( .A1(n688), .A2(n5821), .ZN(n2093) );
  OAI21_X1 U1731 ( .B1(n5506), .B2(n2077), .A(n2094), .ZN(n3533) );
  NAND2_X1 U1732 ( .A1(n689), .A2(n5819), .ZN(n2094) );
  OAI21_X1 U1733 ( .B1(n5503), .B2(n2077), .A(n2095), .ZN(n3532) );
  NAND2_X1 U1734 ( .A1(n690), .A2(n5821), .ZN(n2095) );
  OAI21_X1 U1735 ( .B1(n5500), .B2(n5819), .A(n2096), .ZN(n3531) );
  NAND2_X1 U1736 ( .A1(n691), .A2(n5819), .ZN(n2096) );
  OAI21_X1 U1737 ( .B1(n5497), .B2(n5821), .A(n2097), .ZN(n3530) );
  NAND2_X1 U1738 ( .A1(n692), .A2(n5821), .ZN(n2097) );
  OAI21_X1 U1739 ( .B1(n5494), .B2(n5821), .A(n2098), .ZN(n3529) );
  NAND2_X1 U1740 ( .A1(n693), .A2(n5821), .ZN(n2098) );
  OAI21_X1 U1741 ( .B1(n5491), .B2(n2077), .A(n2099), .ZN(n3528) );
  NAND2_X1 U1742 ( .A1(n694), .A2(n2077), .ZN(n2099) );
  OAI21_X1 U1743 ( .B1(n5488), .B2(n2077), .A(n2100), .ZN(n3527) );
  NAND2_X1 U1744 ( .A1(n695), .A2(n5819), .ZN(n2100) );
  OAI21_X1 U1745 ( .B1(n5485), .B2(n2077), .A(n2101), .ZN(n3526) );
  NAND2_X1 U1746 ( .A1(n696), .A2(n5821), .ZN(n2101) );
  OAI21_X1 U1747 ( .B1(n5482), .B2(n2077), .A(n2102), .ZN(n3525) );
  NAND2_X1 U1748 ( .A1(n697), .A2(n5819), .ZN(n2102) );
  OAI21_X1 U1749 ( .B1(n6082), .B2(n2077), .A(n2103), .ZN(n3524) );
  NAND2_X1 U1750 ( .A1(n698), .A2(n5819), .ZN(n2103) );
  OAI21_X1 U1751 ( .B1(n5476), .B2(n2077), .A(n2104), .ZN(n3523) );
  NAND2_X1 U1752 ( .A1(n699), .A2(n5819), .ZN(n2104) );
  OAI21_X1 U1753 ( .B1(n5473), .B2(n2077), .A(n2105), .ZN(n3522) );
  NAND2_X1 U1754 ( .A1(n700), .A2(n5819), .ZN(n2105) );
  OAI21_X1 U1755 ( .B1(n5470), .B2(n2077), .A(n2106), .ZN(n3521) );
  NAND2_X1 U1756 ( .A1(n701), .A2(n5819), .ZN(n2106) );
  OAI21_X1 U1757 ( .B1(n5467), .B2(n2077), .A(n2107), .ZN(n3520) );
  NAND2_X1 U1758 ( .A1(n702), .A2(n5819), .ZN(n2107) );
  OAI21_X1 U1759 ( .B1(n5463), .B2(n2077), .A(n2108), .ZN(n3519) );
  NAND2_X1 U1760 ( .A1(n703), .A2(n5819), .ZN(n2108) );
  OAI21_X1 U1761 ( .B1(n5461), .B2(n5821), .A(n2109), .ZN(n3518) );
  NAND2_X1 U1762 ( .A1(n704), .A2(n5819), .ZN(n2109) );
  NAND2_X1 U1763 ( .A1(n2110), .A2(n1692), .ZN(n2077) );
  OAI21_X1 U1764 ( .B1(n5554), .B2(n5817), .A(n2112), .ZN(n3517) );
  NAND2_X1 U1765 ( .A1(n2111), .A2(n6302), .ZN(n2112) );
  OAI21_X1 U1766 ( .B1(n5551), .B2(n5818), .A(n2113), .ZN(n3516) );
  NAND2_X1 U1767 ( .A1(n2111), .A2(n6301), .ZN(n2113) );
  OAI21_X1 U1768 ( .B1(n5547), .B2(n5817), .A(n2114), .ZN(n3515) );
  NAND2_X1 U1769 ( .A1(n2111), .A2(n6300), .ZN(n2114) );
  OAI21_X1 U1770 ( .B1(n5545), .B2(n5818), .A(n2115), .ZN(n3514) );
  NAND2_X1 U1771 ( .A1(n2111), .A2(n6299), .ZN(n2115) );
  OAI21_X1 U1772 ( .B1(n5542), .B2(n5817), .A(n2116), .ZN(n3513) );
  NAND2_X1 U1773 ( .A1(n2111), .A2(n6298), .ZN(n2116) );
  OAI21_X1 U1774 ( .B1(n5539), .B2(n5818), .A(n2117), .ZN(n3512) );
  NAND2_X1 U1775 ( .A1(n5818), .A2(n6297), .ZN(n2117) );
  OAI21_X1 U1776 ( .B1(n5536), .B2(n5817), .A(n2118), .ZN(n3511) );
  NAND2_X1 U1777 ( .A1(n5818), .A2(n6296), .ZN(n2118) );
  OAI21_X1 U1778 ( .B1(n5533), .B2(n5818), .A(n2119), .ZN(n3510) );
  NAND2_X1 U1779 ( .A1(n5818), .A2(n6295), .ZN(n2119) );
  OAI21_X1 U1780 ( .B1(n5530), .B2(n5817), .A(n2120), .ZN(n3509) );
  NAND2_X1 U1781 ( .A1(n2111), .A2(n6294), .ZN(n2120) );
  OAI21_X1 U1782 ( .B1(n6098), .B2(n5818), .A(n2121), .ZN(n3508) );
  NAND2_X1 U1783 ( .A1(n5817), .A2(n6293), .ZN(n2121) );
  OAI21_X1 U1784 ( .B1(n5524), .B2(n5817), .A(n2122), .ZN(n3507) );
  NAND2_X1 U1785 ( .A1(n2111), .A2(n6292), .ZN(n2122) );
  OAI21_X1 U1786 ( .B1(n5521), .B2(n5817), .A(n2123), .ZN(n3506) );
  NAND2_X1 U1787 ( .A1(n2111), .A2(n6291), .ZN(n2123) );
  OAI21_X1 U1788 ( .B1(n5518), .B2(n5817), .A(n2124), .ZN(n3505) );
  NAND2_X1 U1789 ( .A1(n2111), .A2(n6290), .ZN(n2124) );
  OAI21_X1 U1790 ( .B1(n5515), .B2(n5817), .A(n2125), .ZN(n3504) );
  NAND2_X1 U1791 ( .A1(n2111), .A2(n6289), .ZN(n2125) );
  OAI21_X1 U1792 ( .B1(n5511), .B2(n5817), .A(n2126), .ZN(n3503) );
  NAND2_X1 U1793 ( .A1(n2111), .A2(n6288), .ZN(n2126) );
  OAI21_X1 U1794 ( .B1(n6092), .B2(n5817), .A(n2127), .ZN(n3502) );
  NAND2_X1 U1795 ( .A1(n2111), .A2(n6287), .ZN(n2127) );
  OAI21_X1 U1796 ( .B1(n5506), .B2(n5817), .A(n2128), .ZN(n3501) );
  NAND2_X1 U1797 ( .A1(n2111), .A2(n6286), .ZN(n2128) );
  OAI21_X1 U1798 ( .B1(n5503), .B2(n5817), .A(n2129), .ZN(n3500) );
  NAND2_X1 U1799 ( .A1(n5818), .A2(n6285), .ZN(n2129) );
  OAI21_X1 U1800 ( .B1(n5500), .B2(n5817), .A(n2131), .ZN(n3499) );
  NAND2_X1 U1801 ( .A1(n5817), .A2(n6284), .ZN(n2131) );
  OAI21_X1 U1802 ( .B1(n5497), .B2(n5817), .A(n2132), .ZN(n3498) );
  NAND2_X1 U1803 ( .A1(n5818), .A2(n6283), .ZN(n2132) );
  OAI21_X1 U1804 ( .B1(n5494), .B2(n5817), .A(n2133), .ZN(n3497) );
  NAND2_X1 U1805 ( .A1(n5817), .A2(n6282), .ZN(n2133) );
  OAI21_X1 U1806 ( .B1(n5491), .B2(n5817), .A(n2134), .ZN(n3496) );
  NAND2_X1 U1807 ( .A1(n5817), .A2(n6281), .ZN(n2134) );
  OAI21_X1 U1808 ( .B1(n5488), .B2(n5818), .A(n2136), .ZN(n3495) );
  NAND2_X1 U1809 ( .A1(n2111), .A2(n6280), .ZN(n2136) );
  OAI21_X1 U1810 ( .B1(n5485), .B2(n5818), .A(n2137), .ZN(n3494) );
  NAND2_X1 U1811 ( .A1(n2111), .A2(n6279), .ZN(n2137) );
  OAI21_X1 U1812 ( .B1(n5482), .B2(n5818), .A(n2138), .ZN(n3493) );
  NAND2_X1 U1813 ( .A1(n2111), .A2(n6278), .ZN(n2138) );
  OAI21_X1 U1814 ( .B1(n6082), .B2(n5818), .A(n2139), .ZN(n3492) );
  NAND2_X1 U1815 ( .A1(n2111), .A2(n6277), .ZN(n2139) );
  OAI21_X1 U1816 ( .B1(n5476), .B2(n5818), .A(n2141), .ZN(n3491) );
  NAND2_X1 U1817 ( .A1(n2111), .A2(n6276), .ZN(n2141) );
  OAI21_X1 U1818 ( .B1(n5473), .B2(n5818), .A(n2142), .ZN(n3490) );
  NAND2_X1 U1819 ( .A1(n2111), .A2(n6275), .ZN(n2142) );
  OAI21_X1 U1820 ( .B1(n5470), .B2(n5818), .A(n2143), .ZN(n3489) );
  NAND2_X1 U1821 ( .A1(n2111), .A2(n6274), .ZN(n2143) );
  OAI21_X1 U1822 ( .B1(n5467), .B2(n5818), .A(n2144), .ZN(n3488) );
  NAND2_X1 U1823 ( .A1(n2111), .A2(n6273), .ZN(n2144) );
  OAI21_X1 U1824 ( .B1(n5463), .B2(n5818), .A(n2146), .ZN(n3487) );
  NAND2_X1 U1825 ( .A1(n2111), .A2(n6272), .ZN(n2146) );
  OAI21_X1 U1826 ( .B1(n5461), .B2(n5818), .A(n2147), .ZN(n3486) );
  NAND2_X1 U1827 ( .A1(n2111), .A2(n6271), .ZN(n2147) );
  NAND2_X1 U1828 ( .A1(n1556), .A2(n1521), .ZN(n2111) );
  OAI21_X1 U1829 ( .B1(n5554), .B2(n2148), .A(n2149), .ZN(n3485) );
  NAND2_X1 U1830 ( .A1(n385), .A2(n5807), .ZN(n2149) );
  OAI21_X1 U1831 ( .B1(n5551), .B2(n5809), .A(n2151), .ZN(n3484) );
  NAND2_X1 U1832 ( .A1(n386), .A2(n5807), .ZN(n2151) );
  OAI21_X1 U1833 ( .B1(n5547), .B2(n2148), .A(n2152), .ZN(n3483) );
  NAND2_X1 U1834 ( .A1(n387), .A2(n5807), .ZN(n2152) );
  OAI21_X1 U1835 ( .B1(n5545), .B2(n5807), .A(n2153), .ZN(n3482) );
  NAND2_X1 U1836 ( .A1(n388), .A2(n5807), .ZN(n2153) );
  OAI21_X1 U1837 ( .B1(n5542), .B2(n2148), .A(n2154), .ZN(n3481) );
  NAND2_X1 U1838 ( .A1(n389), .A2(n5807), .ZN(n2154) );
  OAI21_X1 U1839 ( .B1(n5539), .B2(n5809), .A(n2156), .ZN(n3480) );
  NAND2_X1 U1840 ( .A1(n390), .A2(n5809), .ZN(n2156) );
  OAI21_X1 U1841 ( .B1(n5536), .B2(n2148), .A(n2157), .ZN(n3479) );
  NAND2_X1 U1842 ( .A1(n391), .A2(n5809), .ZN(n2157) );
  OAI21_X1 U1843 ( .B1(n5533), .B2(n5807), .A(n2158), .ZN(n3478) );
  NAND2_X1 U1844 ( .A1(n392), .A2(n5809), .ZN(n2158) );
  OAI21_X1 U1845 ( .B1(n5530), .B2(n2148), .A(n2159), .ZN(n3477) );
  NAND2_X1 U1846 ( .A1(n393), .A2(n5809), .ZN(n2159) );
  OAI21_X1 U1847 ( .B1(n6098), .B2(n5807), .A(n2161), .ZN(n3476) );
  NAND2_X1 U1848 ( .A1(n394), .A2(n5809), .ZN(n2161) );
  OAI21_X1 U1849 ( .B1(n5524), .B2(n5809), .A(n2162), .ZN(n3475) );
  NAND2_X1 U1850 ( .A1(n395), .A2(n5809), .ZN(n2162) );
  OAI21_X1 U1851 ( .B1(n5521), .B2(n2148), .A(n2163), .ZN(n3474) );
  NAND2_X1 U1852 ( .A1(n396), .A2(n5809), .ZN(n2163) );
  OAI21_X1 U1853 ( .B1(n5518), .B2(n2148), .A(n2164), .ZN(n3473) );
  NAND2_X1 U1854 ( .A1(n397), .A2(n5809), .ZN(n2164) );
  OAI21_X1 U1855 ( .B1(n5515), .B2(n2148), .A(n2166), .ZN(n3472) );
  NAND2_X1 U1856 ( .A1(n398), .A2(n5809), .ZN(n2166) );
  OAI21_X1 U1857 ( .B1(n5511), .B2(n2148), .A(n2167), .ZN(n3471) );
  NAND2_X1 U1858 ( .A1(n399), .A2(n5809), .ZN(n2167) );
  OAI21_X1 U1859 ( .B1(n6092), .B2(n2148), .A(n2168), .ZN(n3470) );
  NAND2_X1 U1860 ( .A1(n400), .A2(n5809), .ZN(n2168) );
  OAI21_X1 U1861 ( .B1(n5506), .B2(n2148), .A(n2169), .ZN(n3469) );
  NAND2_X1 U1862 ( .A1(n401), .A2(n5807), .ZN(n2169) );
  OAI21_X1 U1863 ( .B1(n5503), .B2(n2148), .A(n2171), .ZN(n3468) );
  NAND2_X1 U1864 ( .A1(n402), .A2(n5809), .ZN(n2171) );
  OAI21_X1 U1865 ( .B1(n5500), .B2(n5807), .A(n2172), .ZN(n3467) );
  NAND2_X1 U1866 ( .A1(n403), .A2(n5807), .ZN(n2172) );
  OAI21_X1 U1867 ( .B1(n5497), .B2(n5809), .A(n2173), .ZN(n3466) );
  NAND2_X1 U1868 ( .A1(n404), .A2(n5809), .ZN(n2173) );
  OAI21_X1 U1869 ( .B1(n5494), .B2(n5809), .A(n2174), .ZN(n3465) );
  NAND2_X1 U1870 ( .A1(n405), .A2(n5809), .ZN(n2174) );
  OAI21_X1 U1871 ( .B1(n5491), .B2(n2148), .A(n2176), .ZN(n3464) );
  NAND2_X1 U1872 ( .A1(n406), .A2(n2148), .ZN(n2176) );
  OAI21_X1 U1873 ( .B1(n5488), .B2(n2148), .A(n2177), .ZN(n3463) );
  NAND2_X1 U1874 ( .A1(n407), .A2(n5807), .ZN(n2177) );
  OAI21_X1 U1875 ( .B1(n5485), .B2(n2148), .A(n2178), .ZN(n3462) );
  NAND2_X1 U1876 ( .A1(n408), .A2(n5809), .ZN(n2178) );
  OAI21_X1 U1877 ( .B1(n5482), .B2(n2148), .A(n2179), .ZN(n3461) );
  NAND2_X1 U1878 ( .A1(n409), .A2(n5807), .ZN(n2179) );
  OAI21_X1 U1879 ( .B1(n6082), .B2(n2148), .A(n2181), .ZN(n3460) );
  NAND2_X1 U1880 ( .A1(n410), .A2(n5807), .ZN(n2181) );
  OAI21_X1 U1881 ( .B1(n5476), .B2(n2148), .A(n2182), .ZN(n3459) );
  NAND2_X1 U1882 ( .A1(n411), .A2(n5807), .ZN(n2182) );
  OAI21_X1 U1883 ( .B1(n5473), .B2(n2148), .A(n2183), .ZN(n3458) );
  NAND2_X1 U1884 ( .A1(n412), .A2(n5807), .ZN(n2183) );
  OAI21_X1 U1885 ( .B1(n5470), .B2(n2148), .A(n2184), .ZN(n3457) );
  NAND2_X1 U1886 ( .A1(n413), .A2(n5807), .ZN(n2184) );
  OAI21_X1 U1887 ( .B1(n5467), .B2(n2148), .A(n2186), .ZN(n3456) );
  NAND2_X1 U1888 ( .A1(n414), .A2(n5807), .ZN(n2186) );
  OAI21_X1 U1889 ( .B1(n5463), .B2(n2148), .A(n2187), .ZN(n3455) );
  NAND2_X1 U1890 ( .A1(n415), .A2(n5807), .ZN(n2187) );
  OAI21_X1 U1891 ( .B1(n5461), .B2(n5809), .A(n2188), .ZN(n3454) );
  NAND2_X1 U1892 ( .A1(n416), .A2(n5807), .ZN(n2188) );
  NAND2_X1 U1893 ( .A1(n1812), .A2(n1556), .ZN(n2148) );
  OAI21_X1 U1894 ( .B1(n5554), .B2(n5806), .A(n2191), .ZN(n3453) );
  NAND2_X1 U1895 ( .A1(n417), .A2(n2189), .ZN(n2191) );
  OAI21_X1 U1896 ( .B1(n5551), .B2(n5805), .A(n2192), .ZN(n3452) );
  NAND2_X1 U1897 ( .A1(n418), .A2(n2189), .ZN(n2192) );
  OAI21_X1 U1898 ( .B1(n5547), .B2(n5806), .A(n2193), .ZN(n3451) );
  NAND2_X1 U1899 ( .A1(n419), .A2(n2189), .ZN(n2193) );
  OAI21_X1 U1900 ( .B1(n5545), .B2(n5805), .A(n2194), .ZN(n3450) );
  NAND2_X1 U1901 ( .A1(n420), .A2(n2189), .ZN(n2194) );
  OAI21_X1 U1902 ( .B1(n5542), .B2(n5806), .A(n2196), .ZN(n3449) );
  NAND2_X1 U1903 ( .A1(n421), .A2(n2189), .ZN(n2196) );
  OAI21_X1 U1904 ( .B1(n5539), .B2(n5805), .A(n2197), .ZN(n3448) );
  NAND2_X1 U1905 ( .A1(n422), .A2(n5806), .ZN(n2197) );
  OAI21_X1 U1906 ( .B1(n5536), .B2(n5806), .A(n2198), .ZN(n3447) );
  NAND2_X1 U1907 ( .A1(n423), .A2(n5806), .ZN(n2198) );
  OAI21_X1 U1908 ( .B1(n5533), .B2(n5805), .A(n2199), .ZN(n3446) );
  NAND2_X1 U1909 ( .A1(n424), .A2(n2189), .ZN(n2199) );
  OAI21_X1 U1910 ( .B1(n5530), .B2(n5806), .A(n2201), .ZN(n3445) );
  NAND2_X1 U1911 ( .A1(n425), .A2(n2189), .ZN(n2201) );
  OAI21_X1 U1912 ( .B1(n6098), .B2(n5805), .A(n2202), .ZN(n3444) );
  NAND2_X1 U1913 ( .A1(n426), .A2(n2189), .ZN(n2202) );
  OAI21_X1 U1914 ( .B1(n5524), .B2(n5806), .A(n2203), .ZN(n3443) );
  NAND2_X1 U1915 ( .A1(n427), .A2(n2189), .ZN(n2203) );
  OAI21_X1 U1916 ( .B1(n5521), .B2(n5805), .A(n2204), .ZN(n3442) );
  NAND2_X1 U1917 ( .A1(n428), .A2(n2189), .ZN(n2204) );
  OAI21_X1 U1918 ( .B1(n5518), .B2(n5805), .A(n2206), .ZN(n3441) );
  NAND2_X1 U1919 ( .A1(n429), .A2(n2189), .ZN(n2206) );
  OAI21_X1 U1920 ( .B1(n5515), .B2(n5805), .A(n2207), .ZN(n3440) );
  NAND2_X1 U1921 ( .A1(n430), .A2(n2189), .ZN(n2207) );
  OAI21_X1 U1922 ( .B1(n5511), .B2(n5805), .A(n2208), .ZN(n3439) );
  NAND2_X1 U1923 ( .A1(n431), .A2(n2189), .ZN(n2208) );
  OAI21_X1 U1924 ( .B1(n6092), .B2(n5805), .A(n2209), .ZN(n3438) );
  NAND2_X1 U1925 ( .A1(n432), .A2(n2189), .ZN(n2209) );
  OAI21_X1 U1926 ( .B1(n5506), .B2(n5805), .A(n2211), .ZN(n3437) );
  NAND2_X1 U1927 ( .A1(n433), .A2(n2189), .ZN(n2211) );
  OAI21_X1 U1928 ( .B1(n5503), .B2(n5805), .A(n2212), .ZN(n3436) );
  NAND2_X1 U1929 ( .A1(n434), .A2(n5805), .ZN(n2212) );
  OAI21_X1 U1930 ( .B1(n5500), .B2(n5805), .A(n2213), .ZN(n3435) );
  NAND2_X1 U1931 ( .A1(n435), .A2(n5805), .ZN(n2213) );
  OAI21_X1 U1932 ( .B1(n5497), .B2(n5805), .A(n2214), .ZN(n3434) );
  NAND2_X1 U1933 ( .A1(n436), .A2(n5806), .ZN(n2214) );
  OAI21_X1 U1934 ( .B1(n5494), .B2(n5805), .A(n2216), .ZN(n3433) );
  NAND2_X1 U1935 ( .A1(n437), .A2(n5806), .ZN(n2216) );
  OAI21_X1 U1936 ( .B1(n5491), .B2(n5805), .A(n2217), .ZN(n3432) );
  NAND2_X1 U1937 ( .A1(n438), .A2(n5805), .ZN(n2217) );
  OAI21_X1 U1938 ( .B1(n5488), .B2(n5806), .A(n2218), .ZN(n3431) );
  NAND2_X1 U1939 ( .A1(n439), .A2(n2189), .ZN(n2218) );
  OAI21_X1 U1940 ( .B1(n5485), .B2(n5806), .A(n2219), .ZN(n3430) );
  NAND2_X1 U1941 ( .A1(n440), .A2(n2189), .ZN(n2219) );
  OAI21_X1 U1942 ( .B1(n5482), .B2(n5806), .A(n2221), .ZN(n3429) );
  NAND2_X1 U1943 ( .A1(n441), .A2(n2189), .ZN(n2221) );
  OAI21_X1 U1944 ( .B1(n6082), .B2(n5806), .A(n2222), .ZN(n3428) );
  NAND2_X1 U1945 ( .A1(n442), .A2(n2189), .ZN(n2222) );
  OAI21_X1 U1946 ( .B1(n5476), .B2(n5806), .A(n2223), .ZN(n3427) );
  NAND2_X1 U1947 ( .A1(n443), .A2(n2189), .ZN(n2223) );
  OAI21_X1 U1948 ( .B1(n5473), .B2(n5806), .A(n2224), .ZN(n3426) );
  NAND2_X1 U1949 ( .A1(n444), .A2(n2189), .ZN(n2224) );
  OAI21_X1 U1950 ( .B1(n5470), .B2(n5806), .A(n2226), .ZN(n3425) );
  NAND2_X1 U1951 ( .A1(n445), .A2(n5806), .ZN(n2226) );
  OAI21_X1 U1952 ( .B1(n5467), .B2(n5806), .A(n2227), .ZN(n3424) );
  NAND2_X1 U1953 ( .A1(n446), .A2(n5805), .ZN(n2227) );
  OAI21_X1 U1954 ( .B1(n5463), .B2(n5806), .A(n2228), .ZN(n3423) );
  NAND2_X1 U1955 ( .A1(n447), .A2(n2189), .ZN(n2228) );
  OAI21_X1 U1956 ( .B1(n5461), .B2(n5806), .A(n2229), .ZN(n3422) );
  NAND2_X1 U1957 ( .A1(n448), .A2(n5805), .ZN(n2229) );
  NAND2_X1 U1958 ( .A1(n1778), .A2(n1556), .ZN(n2189) );
  OAI21_X1 U1959 ( .B1(n5554), .B2(n5800), .A(n2232), .ZN(n3421) );
  NAND2_X1 U1960 ( .A1(n545), .A2(n2231), .ZN(n2232) );
  OAI21_X1 U1961 ( .B1(n5551), .B2(n5799), .A(n2233), .ZN(n3420) );
  NAND2_X1 U1962 ( .A1(n546), .A2(n2231), .ZN(n2233) );
  OAI21_X1 U1963 ( .B1(n5547), .B2(n5800), .A(n2234), .ZN(n3419) );
  NAND2_X1 U1964 ( .A1(n547), .A2(n2231), .ZN(n2234) );
  OAI21_X1 U1965 ( .B1(n5545), .B2(n5799), .A(n2236), .ZN(n3418) );
  NAND2_X1 U1966 ( .A1(n548), .A2(n2231), .ZN(n2236) );
  OAI21_X1 U1967 ( .B1(n5542), .B2(n5800), .A(n2237), .ZN(n3417) );
  NAND2_X1 U1968 ( .A1(n549), .A2(n2231), .ZN(n2237) );
  OAI21_X1 U1969 ( .B1(n5539), .B2(n5799), .A(n2238), .ZN(n3416) );
  NAND2_X1 U1970 ( .A1(n550), .A2(n2231), .ZN(n2238) );
  OAI21_X1 U1971 ( .B1(n5536), .B2(n5800), .A(n2239), .ZN(n3415) );
  NAND2_X1 U1972 ( .A1(n551), .A2(n5800), .ZN(n2239) );
  OAI21_X1 U1973 ( .B1(n5533), .B2(n5799), .A(n2241), .ZN(n3414) );
  NAND2_X1 U1974 ( .A1(n552), .A2(n5799), .ZN(n2241) );
  OAI21_X1 U1975 ( .B1(n5530), .B2(n5800), .A(n2242), .ZN(n3413) );
  NAND2_X1 U1976 ( .A1(n553), .A2(n2231), .ZN(n2242) );
  OAI21_X1 U1977 ( .B1(n6098), .B2(n5799), .A(n2243), .ZN(n3412) );
  NAND2_X1 U1978 ( .A1(n554), .A2(n2231), .ZN(n2243) );
  OAI21_X1 U1979 ( .B1(n5524), .B2(n5800), .A(n2244), .ZN(n3411) );
  NAND2_X1 U1980 ( .A1(n555), .A2(n2231), .ZN(n2244) );
  OAI21_X1 U1981 ( .B1(n5521), .B2(n5799), .A(n2246), .ZN(n3410) );
  NAND2_X1 U1982 ( .A1(n556), .A2(n2231), .ZN(n2246) );
  OAI21_X1 U1983 ( .B1(n5518), .B2(n5799), .A(n2247), .ZN(n3409) );
  NAND2_X1 U1984 ( .A1(n557), .A2(n2231), .ZN(n2247) );
  OAI21_X1 U1985 ( .B1(n5515), .B2(n5799), .A(n2248), .ZN(n3408) );
  NAND2_X1 U1986 ( .A1(n558), .A2(n2231), .ZN(n2248) );
  OAI21_X1 U1987 ( .B1(n5511), .B2(n5799), .A(n2249), .ZN(n3407) );
  NAND2_X1 U1988 ( .A1(n559), .A2(n2231), .ZN(n2249) );
  OAI21_X1 U1989 ( .B1(n5507), .B2(n5799), .A(n2251), .ZN(n3406) );
  NAND2_X1 U1990 ( .A1(n560), .A2(n2231), .ZN(n2251) );
  OAI21_X1 U1991 ( .B1(n6091), .B2(n5799), .A(n2252), .ZN(n3405) );
  NAND2_X1 U1992 ( .A1(n561), .A2(n5800), .ZN(n2252) );
  OAI21_X1 U1993 ( .B1(n6090), .B2(n5799), .A(n2253), .ZN(n3404) );
  NAND2_X1 U1994 ( .A1(n562), .A2(n2231), .ZN(n2253) );
  OAI21_X1 U1995 ( .B1(n6089), .B2(n5799), .A(n2254), .ZN(n3403) );
  NAND2_X1 U1996 ( .A1(n563), .A2(n5799), .ZN(n2254) );
  OAI21_X1 U1997 ( .B1(n6088), .B2(n5799), .A(n2256), .ZN(n3402) );
  NAND2_X1 U1998 ( .A1(n564), .A2(n5799), .ZN(n2256) );
  OAI21_X1 U1999 ( .B1(n6087), .B2(n5799), .A(n2257), .ZN(n3401) );
  NAND2_X1 U2000 ( .A1(n565), .A2(n5800), .ZN(n2257) );
  OAI21_X1 U2001 ( .B1(n6086), .B2(n5799), .A(n2258), .ZN(n3400) );
  NAND2_X1 U2002 ( .A1(n566), .A2(n5800), .ZN(n2258) );
  OAI21_X1 U2003 ( .B1(n6085), .B2(n5800), .A(n2259), .ZN(n3399) );
  NAND2_X1 U2004 ( .A1(n567), .A2(n2231), .ZN(n2259) );
  OAI21_X1 U2005 ( .B1(n6084), .B2(n5800), .A(n2261), .ZN(n3398) );
  NAND2_X1 U2006 ( .A1(n568), .A2(n2231), .ZN(n2261) );
  OAI21_X1 U2007 ( .B1(n6083), .B2(n5800), .A(n2262), .ZN(n3397) );
  NAND2_X1 U2008 ( .A1(n569), .A2(n2231), .ZN(n2262) );
  OAI21_X1 U2009 ( .B1(n5477), .B2(n5800), .A(n2263), .ZN(n3396) );
  NAND2_X1 U2010 ( .A1(n570), .A2(n2231), .ZN(n2263) );
  OAI21_X1 U2011 ( .B1(n6081), .B2(n5800), .A(n2264), .ZN(n3395) );
  NAND2_X1 U2012 ( .A1(n571), .A2(n2231), .ZN(n2264) );
  OAI21_X1 U2013 ( .B1(n6080), .B2(n5800), .A(n2266), .ZN(n3394) );
  NAND2_X1 U2014 ( .A1(n572), .A2(n2231), .ZN(n2266) );
  OAI21_X1 U2015 ( .B1(n6079), .B2(n5800), .A(n2267), .ZN(n3393) );
  NAND2_X1 U2016 ( .A1(n573), .A2(n2231), .ZN(n2267) );
  OAI21_X1 U2017 ( .B1(n6078), .B2(n5800), .A(n2268), .ZN(n3392) );
  NAND2_X1 U2018 ( .A1(n574), .A2(n5800), .ZN(n2268) );
  OAI21_X1 U2019 ( .B1(n6077), .B2(n5800), .A(n2269), .ZN(n3391) );
  NAND2_X1 U2020 ( .A1(n575), .A2(n5799), .ZN(n2269) );
  OAI21_X1 U2021 ( .B1(n6076), .B2(n5800), .A(n2271), .ZN(n3390) );
  NAND2_X1 U2022 ( .A1(n576), .A2(n5799), .ZN(n2271) );
  NAND2_X1 U2023 ( .A1(n2110), .A2(n1556), .ZN(n2231) );
  NOR2_X1 U2024 ( .A1(n2272), .A2(n6065), .ZN(n1556) );
  OR2_X1 U2025 ( .A1(ADD_WR[4]), .A2(n2273), .ZN(n2272) );
  OAI21_X1 U2026 ( .B1(n6107), .B2(n5794), .A(n2275), .ZN(n3389) );
  NAND2_X1 U2027 ( .A1(n449), .A2(n2274), .ZN(n2275) );
  OAI21_X1 U2028 ( .B1(n6106), .B2(n5793), .A(n2276), .ZN(n3388) );
  NAND2_X1 U2029 ( .A1(n450), .A2(n2274), .ZN(n2276) );
  OAI21_X1 U2030 ( .B1(n6105), .B2(n5794), .A(n2277), .ZN(n3387) );
  NAND2_X1 U2031 ( .A1(n451), .A2(n2274), .ZN(n2277) );
  OAI21_X1 U2032 ( .B1(n6104), .B2(n5793), .A(n2278), .ZN(n3386) );
  NAND2_X1 U2033 ( .A1(n452), .A2(n2274), .ZN(n2278) );
  OAI21_X1 U2034 ( .B1(n6103), .B2(n5794), .A(n2279), .ZN(n3385) );
  NAND2_X1 U2035 ( .A1(n453), .A2(n2274), .ZN(n2279) );
  OAI21_X1 U2036 ( .B1(n6102), .B2(n5793), .A(n2280), .ZN(n3384) );
  NAND2_X1 U2037 ( .A1(n454), .A2(n2274), .ZN(n2280) );
  OAI21_X1 U2038 ( .B1(n6101), .B2(n5794), .A(n2281), .ZN(n3383) );
  NAND2_X1 U2039 ( .A1(n455), .A2(n5794), .ZN(n2281) );
  OAI21_X1 U2040 ( .B1(n6100), .B2(n5793), .A(n2282), .ZN(n3382) );
  NAND2_X1 U2041 ( .A1(n456), .A2(n5793), .ZN(n2282) );
  OAI21_X1 U2042 ( .B1(n6099), .B2(n5794), .A(n2283), .ZN(n3381) );
  NAND2_X1 U2043 ( .A1(n457), .A2(n2274), .ZN(n2283) );
  OAI21_X1 U2044 ( .B1(n5525), .B2(n5793), .A(n2284), .ZN(n3380) );
  NAND2_X1 U2045 ( .A1(n458), .A2(n2274), .ZN(n2284) );
  OAI21_X1 U2046 ( .B1(n6097), .B2(n5794), .A(n2285), .ZN(n3379) );
  NAND2_X1 U2047 ( .A1(n459), .A2(n2274), .ZN(n2285) );
  OAI21_X1 U2048 ( .B1(n6096), .B2(n5793), .A(n2286), .ZN(n3378) );
  NAND2_X1 U2049 ( .A1(n460), .A2(n2274), .ZN(n2286) );
  OAI21_X1 U2050 ( .B1(n6095), .B2(n5793), .A(n2287), .ZN(n3377) );
  NAND2_X1 U2051 ( .A1(n461), .A2(n2274), .ZN(n2287) );
  OAI21_X1 U2052 ( .B1(n6094), .B2(n5793), .A(n2288), .ZN(n3376) );
  NAND2_X1 U2053 ( .A1(n462), .A2(n2274), .ZN(n2288) );
  OAI21_X1 U2054 ( .B1(n6093), .B2(n5793), .A(n2289), .ZN(n3375) );
  NAND2_X1 U2055 ( .A1(n463), .A2(n2274), .ZN(n2289) );
  OAI21_X1 U2056 ( .B1(n5507), .B2(n5793), .A(n2290), .ZN(n3374) );
  NAND2_X1 U2057 ( .A1(n464), .A2(n2274), .ZN(n2290) );
  OAI21_X1 U2058 ( .B1(n6091), .B2(n5793), .A(n2291), .ZN(n3373) );
  NAND2_X1 U2059 ( .A1(n465), .A2(n5794), .ZN(n2291) );
  OAI21_X1 U2060 ( .B1(n6090), .B2(n5793), .A(n2292), .ZN(n3372) );
  NAND2_X1 U2061 ( .A1(n466), .A2(n2274), .ZN(n2292) );
  OAI21_X1 U2062 ( .B1(n6089), .B2(n5793), .A(n2293), .ZN(n3371) );
  NAND2_X1 U2063 ( .A1(n467), .A2(n5793), .ZN(n2293) );
  OAI21_X1 U2064 ( .B1(n6088), .B2(n5793), .A(n2294), .ZN(n3370) );
  NAND2_X1 U2065 ( .A1(n468), .A2(n5793), .ZN(n2294) );
  OAI21_X1 U2066 ( .B1(n6087), .B2(n5793), .A(n2295), .ZN(n3369) );
  NAND2_X1 U2067 ( .A1(n469), .A2(n5794), .ZN(n2295) );
  OAI21_X1 U2068 ( .B1(n6086), .B2(n5793), .A(n2296), .ZN(n3368) );
  NAND2_X1 U2069 ( .A1(n470), .A2(n5794), .ZN(n2296) );
  OAI21_X1 U2070 ( .B1(n6085), .B2(n5794), .A(n2297), .ZN(n3367) );
  NAND2_X1 U2071 ( .A1(n471), .A2(n2274), .ZN(n2297) );
  OAI21_X1 U2072 ( .B1(n6084), .B2(n5794), .A(n2298), .ZN(n3366) );
  NAND2_X1 U2073 ( .A1(n472), .A2(n2274), .ZN(n2298) );
  OAI21_X1 U2074 ( .B1(n6083), .B2(n5794), .A(n2299), .ZN(n3365) );
  NAND2_X1 U2075 ( .A1(n473), .A2(n2274), .ZN(n2299) );
  OAI21_X1 U2076 ( .B1(n5477), .B2(n5794), .A(n2300), .ZN(n3364) );
  NAND2_X1 U2077 ( .A1(n474), .A2(n2274), .ZN(n2300) );
  OAI21_X1 U2078 ( .B1(n6081), .B2(n5794), .A(n2301), .ZN(n3363) );
  NAND2_X1 U2079 ( .A1(n475), .A2(n2274), .ZN(n2301) );
  OAI21_X1 U2080 ( .B1(n6080), .B2(n5794), .A(n2302), .ZN(n3362) );
  NAND2_X1 U2081 ( .A1(n476), .A2(n2274), .ZN(n2302) );
  OAI21_X1 U2082 ( .B1(n6079), .B2(n5794), .A(n2303), .ZN(n3361) );
  NAND2_X1 U2083 ( .A1(n477), .A2(n2274), .ZN(n2303) );
  OAI21_X1 U2084 ( .B1(n6078), .B2(n5794), .A(n2304), .ZN(n3360) );
  NAND2_X1 U2085 ( .A1(n478), .A2(n5794), .ZN(n2304) );
  OAI21_X1 U2086 ( .B1(n6077), .B2(n5794), .A(n2305), .ZN(n3359) );
  NAND2_X1 U2087 ( .A1(n479), .A2(n5793), .ZN(n2305) );
  OAI21_X1 U2088 ( .B1(n6076), .B2(n5794), .A(n2306), .ZN(n3358) );
  NAND2_X1 U2089 ( .A1(n480), .A2(n5793), .ZN(n2306) );
  NAND2_X1 U2090 ( .A1(n1658), .A2(n1520), .ZN(n2274) );
  NOR2_X1 U2092 ( .A1(n6067), .A2(n6066), .ZN(n2307) );
  OAI21_X1 U2093 ( .B1(n6107), .B2(n5785), .A(n2309), .ZN(n3357) );
  NAND2_X1 U2094 ( .A1(n5783), .A2(n6235), .ZN(n2309) );
  OAI21_X1 U2095 ( .B1(n6106), .B2(n5785), .A(n2310), .ZN(n3356) );
  NAND2_X1 U2096 ( .A1(n5783), .A2(n6234), .ZN(n2310) );
  OAI21_X1 U2097 ( .B1(n6105), .B2(n2308), .A(n2311), .ZN(n3355) );
  NAND2_X1 U2098 ( .A1(n5783), .A2(n6233), .ZN(n2311) );
  OAI21_X1 U2099 ( .B1(n6104), .B2(n5783), .A(n2312), .ZN(n3354) );
  NAND2_X1 U2100 ( .A1(n5783), .A2(n6232), .ZN(n2312) );
  OAI21_X1 U2101 ( .B1(n6103), .B2(n2308), .A(n2313), .ZN(n3353) );
  NAND2_X1 U2102 ( .A1(n5783), .A2(n6231), .ZN(n2313) );
  OAI21_X1 U2103 ( .B1(n6102), .B2(n5785), .A(n2314), .ZN(n3352) );
  NAND2_X1 U2104 ( .A1(n5785), .A2(n6230), .ZN(n2314) );
  OAI21_X1 U2105 ( .B1(n6101), .B2(n2308), .A(n2315), .ZN(n3351) );
  NAND2_X1 U2106 ( .A1(n5785), .A2(n6229), .ZN(n2315) );
  OAI21_X1 U2107 ( .B1(n6100), .B2(n2308), .A(n2316), .ZN(n3350) );
  NAND2_X1 U2108 ( .A1(n5785), .A2(n6228), .ZN(n2316) );
  OAI21_X1 U2109 ( .B1(n6099), .B2(n2308), .A(n2317), .ZN(n3349) );
  NAND2_X1 U2110 ( .A1(n5785), .A2(n6227), .ZN(n2317) );
  OAI21_X1 U2111 ( .B1(n5525), .B2(n2308), .A(n2318), .ZN(n3348) );
  NAND2_X1 U2112 ( .A1(n5785), .A2(n6226), .ZN(n2318) );
  OAI21_X1 U2113 ( .B1(n6097), .B2(n2308), .A(n2319), .ZN(n3347) );
  NAND2_X1 U2114 ( .A1(n5785), .A2(n6225), .ZN(n2319) );
  OAI21_X1 U2115 ( .B1(n6096), .B2(n2308), .A(n2320), .ZN(n3346) );
  NAND2_X1 U2116 ( .A1(n5785), .A2(n6224), .ZN(n2320) );
  OAI21_X1 U2117 ( .B1(n6095), .B2(n2308), .A(n2321), .ZN(n3345) );
  NAND2_X1 U2118 ( .A1(n5785), .A2(n6223), .ZN(n2321) );
  OAI21_X1 U2119 ( .B1(n6094), .B2(n2308), .A(n2322), .ZN(n3344) );
  NAND2_X1 U2120 ( .A1(n5785), .A2(n6222), .ZN(n2322) );
  OAI21_X1 U2121 ( .B1(n6093), .B2(n2308), .A(n2323), .ZN(n3343) );
  NAND2_X1 U2122 ( .A1(n5785), .A2(n6221), .ZN(n2323) );
  OAI21_X1 U2123 ( .B1(n5507), .B2(n2308), .A(n2324), .ZN(n3342) );
  NAND2_X1 U2124 ( .A1(n5785), .A2(n6220), .ZN(n2324) );
  OAI21_X1 U2125 ( .B1(n6091), .B2(n5785), .A(n2325), .ZN(n3341) );
  NAND2_X1 U2126 ( .A1(n5783), .A2(n6219), .ZN(n2325) );
  OAI21_X1 U2127 ( .B1(n6090), .B2(n5783), .A(n2326), .ZN(n3340) );
  NAND2_X1 U2128 ( .A1(n5785), .A2(n6218), .ZN(n2326) );
  OAI21_X1 U2129 ( .B1(n6089), .B2(n5785), .A(n2327), .ZN(n3339) );
  NAND2_X1 U2130 ( .A1(n5783), .A2(n6217), .ZN(n2327) );
  OAI21_X1 U2131 ( .B1(n6088), .B2(n2308), .A(n2328), .ZN(n3338) );
  NAND2_X1 U2132 ( .A1(n5785), .A2(n6216), .ZN(n2328) );
  OAI21_X1 U2133 ( .B1(n6087), .B2(n5783), .A(n2329), .ZN(n3337) );
  NAND2_X1 U2134 ( .A1(n5785), .A2(n6215), .ZN(n2329) );
  OAI21_X1 U2135 ( .B1(n6086), .B2(n5783), .A(n2330), .ZN(n3336) );
  NAND2_X1 U2136 ( .A1(n2308), .A2(n6214), .ZN(n2330) );
  OAI21_X1 U2137 ( .B1(n6085), .B2(n2308), .A(n2331), .ZN(n3335) );
  NAND2_X1 U2138 ( .A1(n5783), .A2(n6213), .ZN(n2331) );
  OAI21_X1 U2139 ( .B1(n6084), .B2(n2308), .A(n2332), .ZN(n3334) );
  NAND2_X1 U2140 ( .A1(n5785), .A2(n6212), .ZN(n2332) );
  OAI21_X1 U2141 ( .B1(n6083), .B2(n2308), .A(n2333), .ZN(n3333) );
  NAND2_X1 U2142 ( .A1(n5783), .A2(n6211), .ZN(n2333) );
  OAI21_X1 U2143 ( .B1(n5477), .B2(n2308), .A(n2334), .ZN(n3332) );
  NAND2_X1 U2144 ( .A1(n5783), .A2(n6210), .ZN(n2334) );
  OAI21_X1 U2145 ( .B1(n6081), .B2(n2308), .A(n2335), .ZN(n3331) );
  NAND2_X1 U2146 ( .A1(n5783), .A2(n6209), .ZN(n2335) );
  OAI21_X1 U2147 ( .B1(n6080), .B2(n2308), .A(n2336), .ZN(n3330) );
  NAND2_X1 U2148 ( .A1(n5783), .A2(n6208), .ZN(n2336) );
  OAI21_X1 U2149 ( .B1(n6079), .B2(n2308), .A(n2337), .ZN(n3329) );
  NAND2_X1 U2150 ( .A1(n5783), .A2(n6207), .ZN(n2337) );
  OAI21_X1 U2151 ( .B1(n6078), .B2(n2308), .A(n2338), .ZN(n3328) );
  NAND2_X1 U2152 ( .A1(n5783), .A2(n6206), .ZN(n2338) );
  OAI21_X1 U2153 ( .B1(n6077), .B2(n2308), .A(n2339), .ZN(n3327) );
  NAND2_X1 U2154 ( .A1(n5783), .A2(n6205), .ZN(n2339) );
  OAI21_X1 U2155 ( .B1(n6076), .B2(n5785), .A(n2340), .ZN(n3326) );
  NAND2_X1 U2156 ( .A1(n5783), .A2(n6204), .ZN(n2340) );
  NAND2_X1 U2157 ( .A1(n1624), .A2(n1520), .ZN(n2308) );
  NOR2_X1 U2159 ( .A1(ADD_WR[0]), .A2(n6066), .ZN(n2341) );
  OAI21_X1 U2160 ( .B1(n6107), .B2(n5782), .A(n2343), .ZN(n3325) );
  NAND2_X1 U2161 ( .A1(n577), .A2(n2342), .ZN(n2343) );
  OAI21_X1 U2162 ( .B1(n6106), .B2(n5781), .A(n2344), .ZN(n3324) );
  NAND2_X1 U2163 ( .A1(n578), .A2(n2342), .ZN(n2344) );
  OAI21_X1 U2164 ( .B1(n6105), .B2(n5782), .A(n2345), .ZN(n3323) );
  NAND2_X1 U2165 ( .A1(n579), .A2(n2342), .ZN(n2345) );
  OAI21_X1 U2166 ( .B1(n6104), .B2(n5781), .A(n2346), .ZN(n3322) );
  NAND2_X1 U2167 ( .A1(n580), .A2(n2342), .ZN(n2346) );
  OAI21_X1 U2168 ( .B1(n6103), .B2(n5782), .A(n2347), .ZN(n3321) );
  NAND2_X1 U2169 ( .A1(n581), .A2(n2342), .ZN(n2347) );
  OAI21_X1 U2170 ( .B1(n6102), .B2(n5781), .A(n2348), .ZN(n3320) );
  NAND2_X1 U2171 ( .A1(n582), .A2(n2342), .ZN(n2348) );
  OAI21_X1 U2172 ( .B1(n6101), .B2(n5782), .A(n2349), .ZN(n3319) );
  NAND2_X1 U2173 ( .A1(n583), .A2(n5782), .ZN(n2349) );
  OAI21_X1 U2174 ( .B1(n6100), .B2(n5781), .A(n2350), .ZN(n3318) );
  NAND2_X1 U2175 ( .A1(n584), .A2(n5781), .ZN(n2350) );
  OAI21_X1 U2176 ( .B1(n6099), .B2(n5782), .A(n2351), .ZN(n3317) );
  NAND2_X1 U2177 ( .A1(n585), .A2(n2342), .ZN(n2351) );
  OAI21_X1 U2178 ( .B1(n5525), .B2(n5781), .A(n2353), .ZN(n3316) );
  NAND2_X1 U2179 ( .A1(n586), .A2(n2342), .ZN(n2353) );
  OAI21_X1 U2180 ( .B1(n6097), .B2(n5782), .A(n2354), .ZN(n3315) );
  NAND2_X1 U2181 ( .A1(n587), .A2(n2342), .ZN(n2354) );
  OAI21_X1 U2182 ( .B1(n6096), .B2(n5781), .A(n2356), .ZN(n3314) );
  NAND2_X1 U2183 ( .A1(n588), .A2(n2342), .ZN(n2356) );
  OAI21_X1 U2184 ( .B1(n6095), .B2(n5781), .A(n2357), .ZN(n3313) );
  NAND2_X1 U2185 ( .A1(n589), .A2(n2342), .ZN(n2357) );
  OAI21_X1 U2186 ( .B1(n6094), .B2(n5781), .A(n2359), .ZN(n3312) );
  NAND2_X1 U2187 ( .A1(n590), .A2(n2342), .ZN(n2359) );
  OAI21_X1 U2188 ( .B1(n6093), .B2(n5781), .A(n2360), .ZN(n3311) );
  NAND2_X1 U2189 ( .A1(n591), .A2(n2342), .ZN(n2360) );
  OAI21_X1 U2190 ( .B1(n5507), .B2(n5781), .A(n2362), .ZN(n3310) );
  NAND2_X1 U2191 ( .A1(n592), .A2(n2342), .ZN(n2362) );
  OAI21_X1 U2192 ( .B1(n6091), .B2(n5781), .A(n2363), .ZN(n3309) );
  NAND2_X1 U2193 ( .A1(n593), .A2(n5782), .ZN(n2363) );
  OAI21_X1 U2194 ( .B1(n6090), .B2(n5781), .A(n2365), .ZN(n3308) );
  NAND2_X1 U2195 ( .A1(n594), .A2(n2342), .ZN(n2365) );
  OAI21_X1 U2196 ( .B1(n6089), .B2(n5781), .A(n2366), .ZN(n3307) );
  NAND2_X1 U2197 ( .A1(n595), .A2(n5781), .ZN(n2366) );
  OAI21_X1 U2198 ( .B1(n6088), .B2(n5781), .A(n2368), .ZN(n3306) );
  NAND2_X1 U2199 ( .A1(n596), .A2(n5781), .ZN(n2368) );
  OAI21_X1 U2200 ( .B1(n6087), .B2(n5781), .A(n2369), .ZN(n3305) );
  NAND2_X1 U2201 ( .A1(n597), .A2(n5782), .ZN(n2369) );
  OAI21_X1 U2202 ( .B1(n6086), .B2(n5781), .A(n2371), .ZN(n3304) );
  NAND2_X1 U2203 ( .A1(n598), .A2(n5782), .ZN(n2371) );
  OAI21_X1 U2204 ( .B1(n6085), .B2(n5782), .A(n2372), .ZN(n3303) );
  NAND2_X1 U2205 ( .A1(n599), .A2(n2342), .ZN(n2372) );
  OAI21_X1 U2206 ( .B1(n6084), .B2(n5782), .A(n2374), .ZN(n3302) );
  NAND2_X1 U2207 ( .A1(n600), .A2(n2342), .ZN(n2374) );
  OAI21_X1 U2208 ( .B1(n6083), .B2(n5782), .A(n2375), .ZN(n3301) );
  NAND2_X1 U2209 ( .A1(n601), .A2(n2342), .ZN(n2375) );
  OAI21_X1 U2210 ( .B1(n5477), .B2(n5782), .A(n2377), .ZN(n3300) );
  NAND2_X1 U2211 ( .A1(n602), .A2(n2342), .ZN(n2377) );
  OAI21_X1 U2212 ( .B1(n6081), .B2(n5782), .A(n2378), .ZN(n3299) );
  NAND2_X1 U2213 ( .A1(n603), .A2(n2342), .ZN(n2378) );
  OAI21_X1 U2214 ( .B1(n6080), .B2(n5782), .A(n2380), .ZN(n3298) );
  NAND2_X1 U2215 ( .A1(n604), .A2(n2342), .ZN(n2380) );
  OAI21_X1 U2216 ( .B1(n6079), .B2(n5782), .A(n2381), .ZN(n3297) );
  NAND2_X1 U2217 ( .A1(n605), .A2(n2342), .ZN(n2381) );
  OAI21_X1 U2218 ( .B1(n6078), .B2(n5782), .A(n2383), .ZN(n3296) );
  NAND2_X1 U2219 ( .A1(n606), .A2(n5782), .ZN(n2383) );
  OAI21_X1 U2220 ( .B1(n6077), .B2(n5782), .A(n2384), .ZN(n3295) );
  NAND2_X1 U2221 ( .A1(n607), .A2(n5781), .ZN(n2384) );
  OAI21_X1 U2222 ( .B1(n6076), .B2(n5782), .A(n2385), .ZN(n3294) );
  NAND2_X1 U2223 ( .A1(n608), .A2(n5781), .ZN(n2385) );
  NAND2_X1 U2224 ( .A1(n1590), .A2(n1520), .ZN(n2342) );
  OAI21_X1 U2225 ( .B1(n6107), .B2(n5775), .A(n2387), .ZN(n3293) );
  NAND2_X1 U2226 ( .A1(n2386), .A2(n6139), .ZN(n2387) );
  OAI21_X1 U2227 ( .B1(n6106), .B2(n5776), .A(n2388), .ZN(n3292) );
  NAND2_X1 U2228 ( .A1(n2386), .A2(n6138), .ZN(n2388) );
  OAI21_X1 U2229 ( .B1(n6105), .B2(n5775), .A(n2389), .ZN(n3291) );
  NAND2_X1 U2230 ( .A1(n2386), .A2(n6137), .ZN(n2389) );
  OAI21_X1 U2231 ( .B1(n6104), .B2(n5776), .A(n2390), .ZN(n3290) );
  NAND2_X1 U2232 ( .A1(n2386), .A2(n6136), .ZN(n2390) );
  OAI21_X1 U2233 ( .B1(n6103), .B2(n5775), .A(n2391), .ZN(n3289) );
  NAND2_X1 U2234 ( .A1(n2386), .A2(n6135), .ZN(n2391) );
  OAI21_X1 U2235 ( .B1(n6102), .B2(n5776), .A(n2392), .ZN(n3288) );
  NAND2_X1 U2236 ( .A1(n2386), .A2(n6134), .ZN(n2392) );
  OAI21_X1 U2237 ( .B1(n6101), .B2(n5775), .A(n2393), .ZN(n3287) );
  NAND2_X1 U2238 ( .A1(n5775), .A2(n6133), .ZN(n2393) );
  OAI21_X1 U2239 ( .B1(n6100), .B2(n5776), .A(n2394), .ZN(n3286) );
  NAND2_X1 U2240 ( .A1(n5775), .A2(n6132), .ZN(n2394) );
  OAI21_X1 U2241 ( .B1(n6099), .B2(n5775), .A(n2395), .ZN(n3285) );
  NAND2_X1 U2242 ( .A1(n5776), .A2(n6131), .ZN(n2395) );
  OAI21_X1 U2243 ( .B1(n5525), .B2(n5776), .A(n2396), .ZN(n3284) );
  NAND2_X1 U2244 ( .A1(n2386), .A2(n6130), .ZN(n2396) );
  OAI21_X1 U2245 ( .B1(n6097), .B2(n5775), .A(n2397), .ZN(n3283) );
  NAND2_X1 U2246 ( .A1(n5775), .A2(n6129), .ZN(n2397) );
  OAI21_X1 U2247 ( .B1(n6096), .B2(n5775), .A(n2398), .ZN(n3282) );
  NAND2_X1 U2248 ( .A1(n2386), .A2(n6128), .ZN(n2398) );
  OAI21_X1 U2249 ( .B1(n6095), .B2(n5775), .A(n2399), .ZN(n3281) );
  NAND2_X1 U2250 ( .A1(n2386), .A2(n6127), .ZN(n2399) );
  OAI21_X1 U2251 ( .B1(n6094), .B2(n5775), .A(n2400), .ZN(n3280) );
  NAND2_X1 U2252 ( .A1(n2386), .A2(n6126), .ZN(n2400) );
  OAI21_X1 U2253 ( .B1(n6093), .B2(n5775), .A(n2401), .ZN(n3279) );
  NAND2_X1 U2254 ( .A1(n2386), .A2(n6125), .ZN(n2401) );
  OAI21_X1 U2255 ( .B1(n5507), .B2(n5775), .A(n2402), .ZN(n3278) );
  NAND2_X1 U2256 ( .A1(n2386), .A2(n6124), .ZN(n2402) );
  OAI21_X1 U2257 ( .B1(n6091), .B2(n5775), .A(n2403), .ZN(n3277) );
  NAND2_X1 U2258 ( .A1(n5776), .A2(n6123), .ZN(n2403) );
  OAI21_X1 U2259 ( .B1(n6090), .B2(n5775), .A(n2404), .ZN(n3276) );
  NAND2_X1 U2260 ( .A1(n2386), .A2(n6122), .ZN(n2404) );
  OAI21_X1 U2261 ( .B1(n6089), .B2(n5775), .A(n2405), .ZN(n3275) );
  NAND2_X1 U2262 ( .A1(n5776), .A2(n6121), .ZN(n2405) );
  OAI21_X1 U2263 ( .B1(n6088), .B2(n5775), .A(n2406), .ZN(n3274) );
  NAND2_X1 U2264 ( .A1(n5775), .A2(n6120), .ZN(n2406) );
  OAI21_X1 U2265 ( .B1(n6087), .B2(n5775), .A(n2407), .ZN(n3273) );
  NAND2_X1 U2266 ( .A1(n5776), .A2(n6119), .ZN(n2407) );
  OAI21_X1 U2267 ( .B1(n6086), .B2(n5775), .A(n2408), .ZN(n3272) );
  NAND2_X1 U2268 ( .A1(n5776), .A2(n6118), .ZN(n2408) );
  OAI21_X1 U2269 ( .B1(n6085), .B2(n5776), .A(n2409), .ZN(n3271) );
  NAND2_X1 U2270 ( .A1(n2386), .A2(n6117), .ZN(n2409) );
  OAI21_X1 U2271 ( .B1(n6084), .B2(n5776), .A(n2410), .ZN(n3270) );
  NAND2_X1 U2272 ( .A1(n2386), .A2(n6116), .ZN(n2410) );
  OAI21_X1 U2273 ( .B1(n6083), .B2(n5776), .A(n2411), .ZN(n3269) );
  NAND2_X1 U2274 ( .A1(n2386), .A2(n6115), .ZN(n2411) );
  OAI21_X1 U2275 ( .B1(n5477), .B2(n5776), .A(n2412), .ZN(n3268) );
  NAND2_X1 U2276 ( .A1(n2386), .A2(n6114), .ZN(n2412) );
  OAI21_X1 U2277 ( .B1(n6081), .B2(n5776), .A(n2413), .ZN(n3267) );
  NAND2_X1 U2278 ( .A1(n2386), .A2(n6113), .ZN(n2413) );
  OAI21_X1 U2279 ( .B1(n6080), .B2(n5776), .A(n2414), .ZN(n3266) );
  NAND2_X1 U2280 ( .A1(n2386), .A2(n6112), .ZN(n2414) );
  OAI21_X1 U2281 ( .B1(n6079), .B2(n5776), .A(n2415), .ZN(n3265) );
  NAND2_X1 U2282 ( .A1(n2386), .A2(n6111), .ZN(n2415) );
  OAI21_X1 U2283 ( .B1(n6078), .B2(n5776), .A(n2416), .ZN(n3264) );
  NAND2_X1 U2284 ( .A1(n2386), .A2(n6110), .ZN(n2416) );
  OAI21_X1 U2285 ( .B1(n6077), .B2(n5776), .A(n2417), .ZN(n3263) );
  NAND2_X1 U2286 ( .A1(n2386), .A2(n6109), .ZN(n2417) );
  OAI21_X1 U2287 ( .B1(n6076), .B2(n5776), .A(n2418), .ZN(n3262) );
  NAND2_X1 U2288 ( .A1(n2386), .A2(n6108), .ZN(n2418) );
  NAND2_X1 U2289 ( .A1(n1555), .A2(n1520), .ZN(n2386) );
  NOR2_X1 U2291 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .ZN(n2419) );
  OAI21_X1 U2292 ( .B1(n6107), .B2(n5770), .A(n2421), .ZN(n3261) );
  NAND2_X1 U2293 ( .A1(n609), .A2(n2420), .ZN(n2421) );
  OAI21_X1 U2294 ( .B1(n6106), .B2(n5769), .A(n2422), .ZN(n3260) );
  NAND2_X1 U2295 ( .A1(n610), .A2(n2420), .ZN(n2422) );
  OAI21_X1 U2296 ( .B1(n6105), .B2(n5770), .A(n2423), .ZN(n3259) );
  NAND2_X1 U2297 ( .A1(n611), .A2(n2420), .ZN(n2423) );
  OAI21_X1 U2298 ( .B1(n6104), .B2(n5769), .A(n2424), .ZN(n3258) );
  NAND2_X1 U2299 ( .A1(n612), .A2(n2420), .ZN(n2424) );
  OAI21_X1 U2300 ( .B1(n6103), .B2(n5770), .A(n2425), .ZN(n3257) );
  NAND2_X1 U2301 ( .A1(n613), .A2(n2420), .ZN(n2425) );
  OAI21_X1 U2302 ( .B1(n6102), .B2(n5769), .A(n2426), .ZN(n3256) );
  NAND2_X1 U2303 ( .A1(n614), .A2(n2420), .ZN(n2426) );
  OAI21_X1 U2304 ( .B1(n6101), .B2(n5770), .A(n2427), .ZN(n3255) );
  NAND2_X1 U2305 ( .A1(n615), .A2(n5770), .ZN(n2427) );
  OAI21_X1 U2306 ( .B1(n6100), .B2(n5769), .A(n2428), .ZN(n3254) );
  NAND2_X1 U2307 ( .A1(n616), .A2(n5769), .ZN(n2428) );
  OAI21_X1 U2308 ( .B1(n6099), .B2(n5770), .A(n2429), .ZN(n3253) );
  NAND2_X1 U2309 ( .A1(n617), .A2(n2420), .ZN(n2429) );
  OAI21_X1 U2310 ( .B1(n5525), .B2(n5769), .A(n2430), .ZN(n3252) );
  NAND2_X1 U2311 ( .A1(n618), .A2(n2420), .ZN(n2430) );
  OAI21_X1 U2312 ( .B1(n6097), .B2(n5770), .A(n2431), .ZN(n3251) );
  NAND2_X1 U2313 ( .A1(n619), .A2(n2420), .ZN(n2431) );
  OAI21_X1 U2314 ( .B1(n6096), .B2(n5769), .A(n2432), .ZN(n3250) );
  NAND2_X1 U2315 ( .A1(n620), .A2(n2420), .ZN(n2432) );
  OAI21_X1 U2316 ( .B1(n6095), .B2(n5769), .A(n2433), .ZN(n3249) );
  NAND2_X1 U2317 ( .A1(n621), .A2(n2420), .ZN(n2433) );
  OAI21_X1 U2318 ( .B1(n6094), .B2(n5769), .A(n2434), .ZN(n3248) );
  NAND2_X1 U2319 ( .A1(n622), .A2(n2420), .ZN(n2434) );
  OAI21_X1 U2320 ( .B1(n6093), .B2(n5769), .A(n2435), .ZN(n3247) );
  NAND2_X1 U2321 ( .A1(n623), .A2(n2420), .ZN(n2435) );
  OAI21_X1 U2322 ( .B1(n5507), .B2(n5769), .A(n2436), .ZN(n3246) );
  NAND2_X1 U2323 ( .A1(n624), .A2(n2420), .ZN(n2436) );
  OAI21_X1 U2324 ( .B1(n6091), .B2(n5769), .A(n2437), .ZN(n3245) );
  NAND2_X1 U2325 ( .A1(n625), .A2(n5770), .ZN(n2437) );
  OAI21_X1 U2326 ( .B1(n6090), .B2(n5769), .A(n2438), .ZN(n3244) );
  NAND2_X1 U2327 ( .A1(n626), .A2(n2420), .ZN(n2438) );
  OAI21_X1 U2328 ( .B1(n6089), .B2(n5769), .A(n2439), .ZN(n3243) );
  NAND2_X1 U2329 ( .A1(n627), .A2(n5769), .ZN(n2439) );
  OAI21_X1 U2330 ( .B1(n6088), .B2(n5769), .A(n2440), .ZN(n3242) );
  NAND2_X1 U2331 ( .A1(n628), .A2(n5769), .ZN(n2440) );
  OAI21_X1 U2332 ( .B1(n6087), .B2(n5769), .A(n2441), .ZN(n3241) );
  NAND2_X1 U2333 ( .A1(n629), .A2(n5770), .ZN(n2441) );
  OAI21_X1 U2334 ( .B1(n6086), .B2(n5769), .A(n2442), .ZN(n3240) );
  NAND2_X1 U2335 ( .A1(n630), .A2(n5770), .ZN(n2442) );
  OAI21_X1 U2336 ( .B1(n6085), .B2(n5770), .A(n2443), .ZN(n3239) );
  NAND2_X1 U2337 ( .A1(n631), .A2(n2420), .ZN(n2443) );
  OAI21_X1 U2338 ( .B1(n6084), .B2(n5770), .A(n2444), .ZN(n3238) );
  NAND2_X1 U2339 ( .A1(n632), .A2(n2420), .ZN(n2444) );
  OAI21_X1 U2340 ( .B1(n6083), .B2(n5770), .A(n2445), .ZN(n3237) );
  NAND2_X1 U2341 ( .A1(n633), .A2(n2420), .ZN(n2445) );
  OAI21_X1 U2342 ( .B1(n5477), .B2(n5770), .A(n2446), .ZN(n3236) );
  NAND2_X1 U2343 ( .A1(n634), .A2(n2420), .ZN(n2446) );
  OAI21_X1 U2344 ( .B1(n6081), .B2(n5770), .A(n2447), .ZN(n3235) );
  NAND2_X1 U2345 ( .A1(n635), .A2(n2420), .ZN(n2447) );
  OAI21_X1 U2346 ( .B1(n6080), .B2(n5770), .A(n2448), .ZN(n3234) );
  NAND2_X1 U2347 ( .A1(n636), .A2(n2420), .ZN(n2448) );
  OAI21_X1 U2348 ( .B1(n6079), .B2(n5770), .A(n2449), .ZN(n3233) );
  NAND2_X1 U2349 ( .A1(n637), .A2(n2420), .ZN(n2449) );
  OAI21_X1 U2350 ( .B1(n6078), .B2(n5770), .A(n2450), .ZN(n3232) );
  NAND2_X1 U2351 ( .A1(n638), .A2(n5770), .ZN(n2450) );
  OAI21_X1 U2352 ( .B1(n6077), .B2(n5770), .A(n2451), .ZN(n3231) );
  NAND2_X1 U2353 ( .A1(n639), .A2(n5769), .ZN(n2451) );
  OAI21_X1 U2354 ( .B1(n6076), .B2(n5770), .A(n2452), .ZN(n3230) );
  NAND2_X1 U2355 ( .A1(n640), .A2(n5769), .ZN(n2452) );
  NAND2_X1 U2356 ( .A1(n1778), .A2(n1520), .ZN(n2420) );
  NOR2_X1 U2357 ( .A1(n2453), .A2(n6067), .ZN(n1778) );
  NAND2_X1 U2358 ( .A1(n2454), .A2(n2455), .ZN(n3229) );
  NOR4_X1 U2359 ( .A1(n2456), .A2(n2457), .A3(n2458), .A4(n2459), .ZN(n2455)
         );
  OAI21_X1 U2360 ( .B1(n1423), .B2(n2460), .A(n2461), .ZN(n2459) );
  NAND2_X1 U2361 ( .A1(n5761), .A2(n6452), .ZN(n2461) );
  OAI21_X1 U2362 ( .B1(n6076), .B2(n5758), .A(n2464), .ZN(n2458) );
  AOI22_X1 U2363 ( .A1(n5755), .A2(n6388), .B1(n5752), .B2(n6420), .ZN(n2464)
         );
  NAND2_X1 U2364 ( .A1(n2467), .A2(n2468), .ZN(n2457) );
  AOI22_X1 U2365 ( .A1(n5749), .A2(n2830), .B1(n5746), .B2(n6516), .ZN(n2468)
         );
  AOI22_X1 U2366 ( .A1(n5743), .A2(n6356), .B1(n5740), .B2(n6239), .ZN(n2467)
         );
  AOI22_X1 U2368 ( .A1(n5735), .A2(n6556), .B1(n5734), .B2(n6303), .ZN(n2476)
         );
  AOI22_X1 U2369 ( .A1(n5731), .A2(n6140), .B1(n5728), .B2(n6588), .ZN(n2475)
         );
  AOI22_X1 U2370 ( .A1(n5725), .A2(n6236), .B1(n5722), .B2(n2382), .ZN(n2474)
         );
  AOI22_X1 U2371 ( .A1(n5717), .A2(n640), .B1(n5716), .B2(n480), .ZN(n2473) );
  NOR4_X1 U2372 ( .A1(n2485), .A2(n2486), .A3(n2487), .A4(n2488), .ZN(n2454)
         );
  NAND2_X1 U2373 ( .A1(n2489), .A2(n2490), .ZN(n2488) );
  AOI22_X1 U2374 ( .A1(n5713), .A2(n416), .B1(n2492), .B2(n6172), .ZN(n2490)
         );
  AOI22_X1 U2375 ( .A1(n5707), .A2(n6271), .B1(n5458), .B2(OUT1[31]), .ZN(
        n2489) );
  NAND2_X1 U2376 ( .A1(n2494), .A2(n2495), .ZN(n2487) );
  AOI22_X1 U2377 ( .A1(n5704), .A2(n448), .B1(n5701), .B2(n6108), .ZN(n2495)
         );
  AOI22_X1 U2378 ( .A1(n5698), .A2(n6204), .B1(n5695), .B2(n576), .ZN(n2494)
         );
  NAND2_X1 U2379 ( .A1(n2500), .A2(n2501), .ZN(n2486) );
  AOI22_X1 U2380 ( .A1(n5691), .A2(n704), .B1(n5689), .B2(n672), .ZN(n2501) );
  AOI22_X1 U2381 ( .A1(n5686), .A2(n736), .B1(n5681), .B2(n608), .ZN(n2500) );
  NAND2_X1 U2382 ( .A1(n2506), .A2(n2507), .ZN(n2485) );
  AOI22_X1 U2383 ( .A1(n5680), .A2(n512), .B1(n5677), .B2(n384), .ZN(n2507) );
  AOI22_X1 U2384 ( .A1(n5674), .A2(n544), .B1(n5671), .B2(n352), .ZN(n2506) );
  NAND2_X1 U2385 ( .A1(n2512), .A2(n2513), .ZN(n3228) );
  NOR4_X1 U2386 ( .A1(n2514), .A2(n2515), .A3(n2516), .A4(n2517), .ZN(n2513)
         );
  OAI21_X1 U2387 ( .B1(n1424), .B2(n2460), .A(n2518), .ZN(n2517) );
  NAND2_X1 U2388 ( .A1(n5761), .A2(n6453), .ZN(n2518) );
  OAI21_X1 U2389 ( .B1(n6077), .B2(n5758), .A(n2519), .ZN(n2516) );
  AOI22_X1 U2390 ( .A1(n5755), .A2(n6389), .B1(n5752), .B2(n6421), .ZN(n2519)
         );
  NAND2_X1 U2391 ( .A1(n2520), .A2(n2521), .ZN(n2515) );
  AOI22_X1 U2392 ( .A1(n5749), .A2(n2829), .B1(n5746), .B2(n6517), .ZN(n2521)
         );
  AOI22_X1 U2393 ( .A1(n5743), .A2(n6357), .B1(n5740), .B2(n6240), .ZN(n2520)
         );
  AOI22_X1 U2395 ( .A1(n5735), .A2(n6557), .B1(n5734), .B2(n6304), .ZN(n2525)
         );
  AOI22_X1 U2396 ( .A1(n5731), .A2(n6141), .B1(n5728), .B2(n6589), .ZN(n2524)
         );
  AOI22_X1 U2397 ( .A1(n5725), .A2(n6237), .B1(n5722), .B2(n2379), .ZN(n2523)
         );
  AOI22_X1 U2398 ( .A1(n5717), .A2(n639), .B1(n5716), .B2(n479), .ZN(n2522) );
  NOR4_X1 U2399 ( .A1(n2526), .A2(n2527), .A3(n2528), .A4(n2529), .ZN(n2512)
         );
  NAND2_X1 U2400 ( .A1(n2530), .A2(n2531), .ZN(n2529) );
  AOI22_X1 U2401 ( .A1(n5713), .A2(n415), .B1(n2492), .B2(n6173), .ZN(n2531)
         );
  AOI22_X1 U2402 ( .A1(n5707), .A2(n6272), .B1(n5458), .B2(OUT1[30]), .ZN(
        n2530) );
  NAND2_X1 U2403 ( .A1(n2532), .A2(n2533), .ZN(n2528) );
  AOI22_X1 U2404 ( .A1(n5704), .A2(n447), .B1(n5701), .B2(n6109), .ZN(n2533)
         );
  AOI22_X1 U2405 ( .A1(n5698), .A2(n6205), .B1(n5695), .B2(n575), .ZN(n2532)
         );
  NAND2_X1 U2406 ( .A1(n2534), .A2(n2535), .ZN(n2527) );
  AOI22_X1 U2407 ( .A1(n2502), .A2(n703), .B1(n5689), .B2(n671), .ZN(n2535) );
  AOI22_X1 U2408 ( .A1(n5686), .A2(n735), .B1(n5681), .B2(n607), .ZN(n2534) );
  NAND2_X1 U2409 ( .A1(n2536), .A2(n2537), .ZN(n2526) );
  AOI22_X1 U2410 ( .A1(n5680), .A2(n511), .B1(n5677), .B2(n383), .ZN(n2537) );
  AOI22_X1 U2411 ( .A1(n5674), .A2(n543), .B1(n5671), .B2(n351), .ZN(n2536) );
  NAND2_X1 U2412 ( .A1(n2538), .A2(n2539), .ZN(n3227) );
  NOR4_X1 U2413 ( .A1(n2540), .A2(n2541), .A3(n2542), .A4(n2543), .ZN(n2539)
         );
  OAI21_X1 U2414 ( .B1(n1425), .B2(n2460), .A(n2544), .ZN(n2543) );
  NAND2_X1 U2415 ( .A1(n5761), .A2(n6454), .ZN(n2544) );
  OAI21_X1 U2416 ( .B1(n6078), .B2(n5758), .A(n2545), .ZN(n2542) );
  AOI22_X1 U2417 ( .A1(n5755), .A2(n6390), .B1(n5752), .B2(n6422), .ZN(n2545)
         );
  NAND2_X1 U2418 ( .A1(n2546), .A2(n2547), .ZN(n2541) );
  AOI22_X1 U2419 ( .A1(n5749), .A2(n2828), .B1(n5746), .B2(n6518), .ZN(n2547)
         );
  AOI22_X1 U2420 ( .A1(n5743), .A2(n6358), .B1(n5740), .B2(n6241), .ZN(n2546)
         );
  AOI22_X1 U2422 ( .A1(n5735), .A2(n6558), .B1(n5734), .B2(n6305), .ZN(n2551)
         );
  AOI22_X1 U2423 ( .A1(n5731), .A2(n6142), .B1(n5728), .B2(n6590), .ZN(n2550)
         );
  AOI22_X1 U2424 ( .A1(n5725), .A2(n6238), .B1(n5722), .B2(n2376), .ZN(n2549)
         );
  AOI22_X1 U2425 ( .A1(n5717), .A2(n638), .B1(n5716), .B2(n478), .ZN(n2548) );
  NOR4_X1 U2426 ( .A1(n2552), .A2(n2553), .A3(n2554), .A4(n2555), .ZN(n2538)
         );
  NAND2_X1 U2427 ( .A1(n2556), .A2(n2557), .ZN(n2555) );
  AOI22_X1 U2428 ( .A1(n5713), .A2(n414), .B1(n2492), .B2(n6174), .ZN(n2557)
         );
  AOI22_X1 U2429 ( .A1(n5707), .A2(n6273), .B1(n5458), .B2(OUT1[29]), .ZN(
        n2556) );
  NAND2_X1 U2430 ( .A1(n2558), .A2(n2559), .ZN(n2554) );
  AOI22_X1 U2431 ( .A1(n5704), .A2(n446), .B1(n5701), .B2(n6110), .ZN(n2559)
         );
  AOI22_X1 U2432 ( .A1(n5698), .A2(n6206), .B1(n5695), .B2(n574), .ZN(n2558)
         );
  NAND2_X1 U2433 ( .A1(n2560), .A2(n2561), .ZN(n2553) );
  AOI22_X1 U2434 ( .A1(n2502), .A2(n702), .B1(n5689), .B2(n670), .ZN(n2561) );
  AOI22_X1 U2435 ( .A1(n5686), .A2(n734), .B1(n5681), .B2(n606), .ZN(n2560) );
  NAND2_X1 U2436 ( .A1(n2562), .A2(n2563), .ZN(n2552) );
  AOI22_X1 U2437 ( .A1(n5680), .A2(n510), .B1(n5677), .B2(n382), .ZN(n2563) );
  AOI22_X1 U2438 ( .A1(n5674), .A2(n542), .B1(n5671), .B2(n350), .ZN(n2562) );
  NAND2_X1 U2439 ( .A1(n2564), .A2(n2565), .ZN(n3226) );
  NOR4_X1 U2440 ( .A1(n2566), .A2(n2567), .A3(n2568), .A4(n2569), .ZN(n2565)
         );
  OAI21_X1 U2441 ( .B1(n1426), .B2(n2460), .A(n2570), .ZN(n2569) );
  NAND2_X1 U2442 ( .A1(n5761), .A2(n6455), .ZN(n2570) );
  OAI21_X1 U2443 ( .B1(n6079), .B2(n5758), .A(n2571), .ZN(n2568) );
  AOI22_X1 U2444 ( .A1(n5755), .A2(n6391), .B1(n5752), .B2(n6423), .ZN(n2571)
         );
  NAND2_X1 U2445 ( .A1(n2572), .A2(n2573), .ZN(n2567) );
  AOI22_X1 U2446 ( .A1(n5749), .A2(n2827), .B1(n5746), .B2(n6519), .ZN(n2573)
         );
  AOI22_X1 U2447 ( .A1(n5743), .A2(n6359), .B1(n5740), .B2(n6242), .ZN(n2572)
         );
  AOI22_X1 U2449 ( .A1(n5735), .A2(n6559), .B1(n5734), .B2(n6306), .ZN(n2577)
         );
  AOI22_X1 U2450 ( .A1(n5731), .A2(n6143), .B1(n5728), .B2(n6591), .ZN(n2576)
         );
  AOI22_X1 U2451 ( .A1(n5725), .A2(n2270), .B1(n5722), .B2(n2373), .ZN(n2575)
         );
  AOI22_X1 U2452 ( .A1(n5717), .A2(n637), .B1(n5716), .B2(n477), .ZN(n2574) );
  NOR4_X1 U2453 ( .A1(n2578), .A2(n2579), .A3(n2580), .A4(n2581), .ZN(n2564)
         );
  NAND2_X1 U2454 ( .A1(n2582), .A2(n2583), .ZN(n2581) );
  AOI22_X1 U2455 ( .A1(n5713), .A2(n413), .B1(n2492), .B2(n6175), .ZN(n2583)
         );
  AOI22_X1 U2456 ( .A1(n5707), .A2(n6274), .B1(n5458), .B2(OUT1[28]), .ZN(
        n2582) );
  NAND2_X1 U2457 ( .A1(n2584), .A2(n2585), .ZN(n2580) );
  AOI22_X1 U2458 ( .A1(n5704), .A2(n445), .B1(n5701), .B2(n6111), .ZN(n2585)
         );
  AOI22_X1 U2459 ( .A1(n5698), .A2(n6207), .B1(n5695), .B2(n573), .ZN(n2584)
         );
  NAND2_X1 U2460 ( .A1(n2586), .A2(n2587), .ZN(n2579) );
  AOI22_X1 U2461 ( .A1(n2502), .A2(n701), .B1(n5689), .B2(n669), .ZN(n2587) );
  AOI22_X1 U2462 ( .A1(n5686), .A2(n733), .B1(n5681), .B2(n605), .ZN(n2586) );
  NAND2_X1 U2463 ( .A1(n2588), .A2(n2589), .ZN(n2578) );
  AOI22_X1 U2464 ( .A1(n5680), .A2(n509), .B1(n5677), .B2(n381), .ZN(n2589) );
  AOI22_X1 U2465 ( .A1(n5674), .A2(n541), .B1(n5671), .B2(n349), .ZN(n2588) );
  NAND2_X1 U2466 ( .A1(n2590), .A2(n2591), .ZN(n3225) );
  NOR4_X1 U2467 ( .A1(n2592), .A2(n2593), .A3(n2594), .A4(n2595), .ZN(n2591)
         );
  OAI21_X1 U2468 ( .B1(n1427), .B2(n2460), .A(n2596), .ZN(n2595) );
  NAND2_X1 U2469 ( .A1(n5761), .A2(n6456), .ZN(n2596) );
  OAI21_X1 U2470 ( .B1(n6080), .B2(n5758), .A(n2597), .ZN(n2594) );
  AOI22_X1 U2471 ( .A1(n5755), .A2(n6392), .B1(n5752), .B2(n6424), .ZN(n2597)
         );
  NAND2_X1 U2472 ( .A1(n2598), .A2(n2599), .ZN(n2593) );
  AOI22_X1 U2473 ( .A1(n5749), .A2(n2826), .B1(n5746), .B2(n6520), .ZN(n2599)
         );
  AOI22_X1 U2474 ( .A1(n5743), .A2(n6360), .B1(n5740), .B2(n6243), .ZN(n2598)
         );
  AOI22_X1 U2476 ( .A1(n5735), .A2(n6560), .B1(n5734), .B2(n6307), .ZN(n2603)
         );
  AOI22_X1 U2477 ( .A1(n5731), .A2(n6144), .B1(n5728), .B2(n6592), .ZN(n2602)
         );
  AOI22_X1 U2478 ( .A1(n5725), .A2(n2265), .B1(n5722), .B2(n2370), .ZN(n2601)
         );
  AOI22_X1 U2479 ( .A1(n5717), .A2(n636), .B1(n5716), .B2(n476), .ZN(n2600) );
  NOR4_X1 U2480 ( .A1(n2604), .A2(n2605), .A3(n2606), .A4(n2607), .ZN(n2590)
         );
  NAND2_X1 U2481 ( .A1(n2608), .A2(n2609), .ZN(n2607) );
  AOI22_X1 U2482 ( .A1(n5713), .A2(n412), .B1(n2492), .B2(n6176), .ZN(n2609)
         );
  AOI22_X1 U2483 ( .A1(n5707), .A2(n6275), .B1(n5458), .B2(OUT1[27]), .ZN(
        n2608) );
  NAND2_X1 U2484 ( .A1(n2610), .A2(n2611), .ZN(n2606) );
  AOI22_X1 U2485 ( .A1(n5704), .A2(n444), .B1(n5701), .B2(n6112), .ZN(n2611)
         );
  AOI22_X1 U2486 ( .A1(n5698), .A2(n6208), .B1(n5695), .B2(n572), .ZN(n2610)
         );
  NAND2_X1 U2487 ( .A1(n2612), .A2(n2613), .ZN(n2605) );
  AOI22_X1 U2488 ( .A1(n2502), .A2(n700), .B1(n5689), .B2(n668), .ZN(n2613) );
  AOI22_X1 U2489 ( .A1(n5686), .A2(n732), .B1(n5681), .B2(n604), .ZN(n2612) );
  NAND2_X1 U2490 ( .A1(n2614), .A2(n2615), .ZN(n2604) );
  AOI22_X1 U2491 ( .A1(n5680), .A2(n508), .B1(n5677), .B2(n380), .ZN(n2615) );
  AOI22_X1 U2492 ( .A1(n5674), .A2(n540), .B1(n5671), .B2(n348), .ZN(n2614) );
  NAND2_X1 U2493 ( .A1(n2616), .A2(n2617), .ZN(n3224) );
  NOR4_X1 U2494 ( .A1(n2618), .A2(n2619), .A3(n2620), .A4(n2621), .ZN(n2617)
         );
  OAI21_X1 U2495 ( .B1(n1428), .B2(n2460), .A(n2622), .ZN(n2621) );
  NAND2_X1 U2496 ( .A1(n5761), .A2(n6457), .ZN(n2622) );
  OAI21_X1 U2497 ( .B1(n6081), .B2(n5758), .A(n2623), .ZN(n2620) );
  AOI22_X1 U2498 ( .A1(n5755), .A2(n6393), .B1(n5752), .B2(n6425), .ZN(n2623)
         );
  NAND2_X1 U2499 ( .A1(n2624), .A2(n2625), .ZN(n2619) );
  AOI22_X1 U2500 ( .A1(n5749), .A2(n2825), .B1(n5746), .B2(n6521), .ZN(n2625)
         );
  AOI22_X1 U2501 ( .A1(n5743), .A2(n6361), .B1(n5740), .B2(n6244), .ZN(n2624)
         );
  AOI22_X1 U2503 ( .A1(n5735), .A2(n6561), .B1(n5734), .B2(n6308), .ZN(n2629)
         );
  AOI22_X1 U2504 ( .A1(n5731), .A2(n6145), .B1(n5728), .B2(n6593), .ZN(n2628)
         );
  AOI22_X1 U2505 ( .A1(n5725), .A2(n2260), .B1(n5722), .B2(n2367), .ZN(n2627)
         );
  AOI22_X1 U2506 ( .A1(n5717), .A2(n635), .B1(n5716), .B2(n475), .ZN(n2626) );
  NOR4_X1 U2507 ( .A1(n2630), .A2(n2631), .A3(n2632), .A4(n2633), .ZN(n2616)
         );
  NAND2_X1 U2508 ( .A1(n2634), .A2(n2635), .ZN(n2633) );
  AOI22_X1 U2509 ( .A1(n5713), .A2(n411), .B1(n2492), .B2(n6177), .ZN(n2635)
         );
  AOI22_X1 U2510 ( .A1(n5707), .A2(n6276), .B1(n5458), .B2(OUT1[26]), .ZN(
        n2634) );
  NAND2_X1 U2511 ( .A1(n2636), .A2(n2637), .ZN(n2632) );
  AOI22_X1 U2512 ( .A1(n5704), .A2(n443), .B1(n5701), .B2(n6113), .ZN(n2637)
         );
  AOI22_X1 U2513 ( .A1(n5698), .A2(n6209), .B1(n5695), .B2(n571), .ZN(n2636)
         );
  NAND2_X1 U2514 ( .A1(n2638), .A2(n2639), .ZN(n2631) );
  AOI22_X1 U2515 ( .A1(n2502), .A2(n699), .B1(n5689), .B2(n667), .ZN(n2639) );
  AOI22_X1 U2516 ( .A1(n5686), .A2(n731), .B1(n5681), .B2(n603), .ZN(n2638) );
  NAND2_X1 U2517 ( .A1(n2640), .A2(n2641), .ZN(n2630) );
  AOI22_X1 U2518 ( .A1(n5680), .A2(n507), .B1(n5677), .B2(n379), .ZN(n2641) );
  AOI22_X1 U2519 ( .A1(n5674), .A2(n539), .B1(n5671), .B2(n347), .ZN(n2640) );
  NAND2_X1 U2520 ( .A1(n2642), .A2(n2643), .ZN(n3223) );
  NOR4_X1 U2521 ( .A1(n2644), .A2(n2645), .A3(n2646), .A4(n2647), .ZN(n2643)
         );
  OAI21_X1 U2522 ( .B1(n1429), .B2(n2460), .A(n2648), .ZN(n2647) );
  NAND2_X1 U2523 ( .A1(n5761), .A2(n6458), .ZN(n2648) );
  OAI21_X1 U2524 ( .B1(n5477), .B2(n5758), .A(n2649), .ZN(n2646) );
  AOI22_X1 U2525 ( .A1(n5755), .A2(n6394), .B1(n5752), .B2(n6426), .ZN(n2649)
         );
  NAND2_X1 U2526 ( .A1(n2650), .A2(n2651), .ZN(n2645) );
  AOI22_X1 U2527 ( .A1(n5749), .A2(n2824), .B1(n5746), .B2(n6522), .ZN(n2651)
         );
  AOI22_X1 U2528 ( .A1(n5743), .A2(n6362), .B1(n5740), .B2(n6245), .ZN(n2650)
         );
  AOI22_X1 U2530 ( .A1(n5735), .A2(n6562), .B1(n5734), .B2(n6309), .ZN(n2655)
         );
  AOI22_X1 U2531 ( .A1(n5731), .A2(n6146), .B1(n5728), .B2(n6594), .ZN(n2654)
         );
  AOI22_X1 U2532 ( .A1(n5725), .A2(n2255), .B1(n5722), .B2(n2364), .ZN(n2653)
         );
  AOI22_X1 U2533 ( .A1(n5717), .A2(n634), .B1(n5716), .B2(n474), .ZN(n2652) );
  NOR4_X1 U2534 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(n2642)
         );
  NAND2_X1 U2535 ( .A1(n2660), .A2(n2661), .ZN(n2659) );
  AOI22_X1 U2536 ( .A1(n5713), .A2(n410), .B1(n2492), .B2(n6178), .ZN(n2661)
         );
  AOI22_X1 U2537 ( .A1(n5707), .A2(n6277), .B1(n5458), .B2(OUT1[25]), .ZN(
        n2660) );
  NAND2_X1 U2538 ( .A1(n2662), .A2(n2663), .ZN(n2658) );
  AOI22_X1 U2539 ( .A1(n5704), .A2(n442), .B1(n5701), .B2(n6114), .ZN(n2663)
         );
  AOI22_X1 U2540 ( .A1(n5698), .A2(n6210), .B1(n5695), .B2(n570), .ZN(n2662)
         );
  NAND2_X1 U2541 ( .A1(n2664), .A2(n2665), .ZN(n2657) );
  AOI22_X1 U2542 ( .A1(n2502), .A2(n698), .B1(n5689), .B2(n666), .ZN(n2665) );
  AOI22_X1 U2543 ( .A1(n5686), .A2(n730), .B1(n5681), .B2(n602), .ZN(n2664) );
  NAND2_X1 U2544 ( .A1(n2666), .A2(n2667), .ZN(n2656) );
  AOI22_X1 U2545 ( .A1(n5680), .A2(n506), .B1(n5677), .B2(n378), .ZN(n2667) );
  AOI22_X1 U2546 ( .A1(n5674), .A2(n538), .B1(n5671), .B2(n346), .ZN(n2666) );
  NAND2_X1 U2547 ( .A1(n2668), .A2(n2669), .ZN(n3222) );
  NOR4_X1 U2548 ( .A1(n2670), .A2(n2671), .A3(n2672), .A4(n2673), .ZN(n2669)
         );
  OAI21_X1 U2549 ( .B1(n1430), .B2(n2460), .A(n2674), .ZN(n2673) );
  NAND2_X1 U2550 ( .A1(n5761), .A2(n6459), .ZN(n2674) );
  OAI21_X1 U2551 ( .B1(n6083), .B2(n5758), .A(n2675), .ZN(n2672) );
  AOI22_X1 U2552 ( .A1(n5755), .A2(n6395), .B1(n5752), .B2(n6427), .ZN(n2675)
         );
  NAND2_X1 U2553 ( .A1(n2676), .A2(n2677), .ZN(n2671) );
  AOI22_X1 U2554 ( .A1(n5749), .A2(n2823), .B1(n5746), .B2(n6523), .ZN(n2677)
         );
  AOI22_X1 U2555 ( .A1(n5743), .A2(n6363), .B1(n5740), .B2(n6246), .ZN(n2676)
         );
  AOI22_X1 U2557 ( .A1(n5735), .A2(n6563), .B1(n5734), .B2(n6310), .ZN(n2681)
         );
  AOI22_X1 U2558 ( .A1(n5731), .A2(n6147), .B1(n5728), .B2(n6595), .ZN(n2680)
         );
  AOI22_X1 U2559 ( .A1(n5725), .A2(n2250), .B1(n5722), .B2(n2361), .ZN(n2679)
         );
  AOI22_X1 U2560 ( .A1(n5717), .A2(n633), .B1(n5716), .B2(n473), .ZN(n2678) );
  NOR4_X1 U2561 ( .A1(n2682), .A2(n2683), .A3(n2684), .A4(n2685), .ZN(n2668)
         );
  NAND2_X1 U2562 ( .A1(n2686), .A2(n2687), .ZN(n2685) );
  AOI22_X1 U2563 ( .A1(n5713), .A2(n409), .B1(n2492), .B2(n6179), .ZN(n2687)
         );
  AOI22_X1 U2564 ( .A1(n5707), .A2(n6278), .B1(n5458), .B2(OUT1[24]), .ZN(
        n2686) );
  NAND2_X1 U2565 ( .A1(n2688), .A2(n2689), .ZN(n2684) );
  AOI22_X1 U2566 ( .A1(n5704), .A2(n441), .B1(n5701), .B2(n6115), .ZN(n2689)
         );
  AOI22_X1 U2567 ( .A1(n5698), .A2(n6211), .B1(n5695), .B2(n569), .ZN(n2688)
         );
  NAND2_X1 U2568 ( .A1(n2690), .A2(n2691), .ZN(n2683) );
  AOI22_X1 U2569 ( .A1(n2502), .A2(n697), .B1(n5689), .B2(n665), .ZN(n2691) );
  AOI22_X1 U2570 ( .A1(n5686), .A2(n729), .B1(n5681), .B2(n601), .ZN(n2690) );
  NAND2_X1 U2571 ( .A1(n2692), .A2(n2693), .ZN(n2682) );
  AOI22_X1 U2572 ( .A1(n5680), .A2(n505), .B1(n5677), .B2(n377), .ZN(n2693) );
  AOI22_X1 U2573 ( .A1(n5674), .A2(n537), .B1(n5671), .B2(n345), .ZN(n2692) );
  NAND2_X1 U2574 ( .A1(n2694), .A2(n2695), .ZN(n3221) );
  NOR4_X1 U2575 ( .A1(n2696), .A2(n2697), .A3(n2698), .A4(n2699), .ZN(n2695)
         );
  OAI21_X1 U2576 ( .B1(n1431), .B2(n2460), .A(n2700), .ZN(n2699) );
  NAND2_X1 U2577 ( .A1(n5761), .A2(n6460), .ZN(n2700) );
  OAI21_X1 U2578 ( .B1(n6084), .B2(n5758), .A(n2701), .ZN(n2698) );
  AOI22_X1 U2579 ( .A1(n5755), .A2(n6396), .B1(n5752), .B2(n6428), .ZN(n2701)
         );
  NAND2_X1 U2580 ( .A1(n2702), .A2(n2703), .ZN(n2697) );
  AOI22_X1 U2581 ( .A1(n5749), .A2(n2822), .B1(n5746), .B2(n6524), .ZN(n2703)
         );
  AOI22_X1 U2582 ( .A1(n5743), .A2(n6364), .B1(n5740), .B2(n6247), .ZN(n2702)
         );
  AOI22_X1 U2584 ( .A1(n5735), .A2(n6564), .B1(n5734), .B2(n6311), .ZN(n2707)
         );
  AOI22_X1 U2585 ( .A1(n5731), .A2(n6148), .B1(n5728), .B2(n6596), .ZN(n2706)
         );
  AOI22_X1 U2586 ( .A1(n5725), .A2(n2245), .B1(n5722), .B2(n2358), .ZN(n2705)
         );
  AOI22_X1 U2587 ( .A1(n2483), .A2(n632), .B1(n5716), .B2(n472), .ZN(n2704) );
  NOR4_X1 U2588 ( .A1(n2708), .A2(n2709), .A3(n2710), .A4(n2711), .ZN(n2694)
         );
  NAND2_X1 U2589 ( .A1(n2712), .A2(n2713), .ZN(n2711) );
  AOI22_X1 U2590 ( .A1(n5713), .A2(n408), .B1(n2492), .B2(n6180), .ZN(n2713)
         );
  AOI22_X1 U2591 ( .A1(n5707), .A2(n6279), .B1(n5458), .B2(OUT1[23]), .ZN(
        n2712) );
  NAND2_X1 U2592 ( .A1(n2714), .A2(n2715), .ZN(n2710) );
  AOI22_X1 U2593 ( .A1(n5704), .A2(n440), .B1(n5701), .B2(n6116), .ZN(n2715)
         );
  AOI22_X1 U2594 ( .A1(n5698), .A2(n6212), .B1(n5695), .B2(n568), .ZN(n2714)
         );
  NAND2_X1 U2595 ( .A1(n2716), .A2(n2717), .ZN(n2709) );
  AOI22_X1 U2596 ( .A1(n2502), .A2(n696), .B1(n5689), .B2(n664), .ZN(n2717) );
  AOI22_X1 U2597 ( .A1(n5686), .A2(n728), .B1(n5681), .B2(n600), .ZN(n2716) );
  NAND2_X1 U2598 ( .A1(n2718), .A2(n2719), .ZN(n2708) );
  AOI22_X1 U2599 ( .A1(n5680), .A2(n504), .B1(n5677), .B2(n376), .ZN(n2719) );
  AOI22_X1 U2600 ( .A1(n5674), .A2(n536), .B1(n5671), .B2(n344), .ZN(n2718) );
  NAND2_X1 U2601 ( .A1(n2720), .A2(n2721), .ZN(n3220) );
  NOR4_X1 U2602 ( .A1(n2722), .A2(n2723), .A3(n2724), .A4(n2725), .ZN(n2721)
         );
  OAI21_X1 U2603 ( .B1(n1432), .B2(n2460), .A(n2726), .ZN(n2725) );
  NAND2_X1 U2604 ( .A1(n5761), .A2(n6461), .ZN(n2726) );
  OAI21_X1 U2605 ( .B1(n6085), .B2(n5758), .A(n2727), .ZN(n2724) );
  AOI22_X1 U2606 ( .A1(n5755), .A2(n6397), .B1(n5752), .B2(n6429), .ZN(n2727)
         );
  NAND2_X1 U2607 ( .A1(n2728), .A2(n2729), .ZN(n2723) );
  AOI22_X1 U2608 ( .A1(n5749), .A2(n2821), .B1(n5746), .B2(n6525), .ZN(n2729)
         );
  AOI22_X1 U2609 ( .A1(n5743), .A2(n6365), .B1(n5740), .B2(n6248), .ZN(n2728)
         );
  AOI22_X1 U2611 ( .A1(n2477), .A2(n6565), .B1(n5734), .B2(n6312), .ZN(n2733)
         );
  AOI22_X1 U2612 ( .A1(n5731), .A2(n6149), .B1(n5728), .B2(n6597), .ZN(n2732)
         );
  AOI22_X1 U2613 ( .A1(n5725), .A2(n2240), .B1(n5722), .B2(n2355), .ZN(n2731)
         );
  AOI22_X1 U2614 ( .A1(n5717), .A2(n631), .B1(n5716), .B2(n471), .ZN(n2730) );
  NOR4_X1 U2615 ( .A1(n2734), .A2(n2735), .A3(n2736), .A4(n2737), .ZN(n2720)
         );
  NAND2_X1 U2616 ( .A1(n2738), .A2(n2739), .ZN(n2737) );
  AOI22_X1 U2617 ( .A1(n5713), .A2(n407), .B1(n2492), .B2(n6181), .ZN(n2739)
         );
  AOI22_X1 U2618 ( .A1(n5707), .A2(n6280), .B1(n5458), .B2(OUT1[22]), .ZN(
        n2738) );
  NAND2_X1 U2619 ( .A1(n2740), .A2(n2741), .ZN(n2736) );
  AOI22_X1 U2620 ( .A1(n5704), .A2(n439), .B1(n5701), .B2(n6117), .ZN(n2741)
         );
  AOI22_X1 U2621 ( .A1(n5698), .A2(n6213), .B1(n5695), .B2(n567), .ZN(n2740)
         );
  NAND2_X1 U2622 ( .A1(n2742), .A2(n2743), .ZN(n2735) );
  AOI22_X1 U2623 ( .A1(n2502), .A2(n695), .B1(n5689), .B2(n663), .ZN(n2743) );
  AOI22_X1 U2624 ( .A1(n5686), .A2(n727), .B1(n5681), .B2(n599), .ZN(n2742) );
  NAND2_X1 U2625 ( .A1(n2744), .A2(n2745), .ZN(n2734) );
  AOI22_X1 U2626 ( .A1(n5680), .A2(n503), .B1(n5677), .B2(n375), .ZN(n2745) );
  AOI22_X1 U2627 ( .A1(n5674), .A2(n535), .B1(n5671), .B2(n343), .ZN(n2744) );
  NAND2_X1 U2628 ( .A1(n2746), .A2(n2747), .ZN(n3219) );
  NOR4_X1 U2629 ( .A1(n2748), .A2(n2749), .A3(n2750), .A4(n2751), .ZN(n2747)
         );
  OAI21_X1 U2630 ( .B1(n1433), .B2(n5763), .A(n2752), .ZN(n2751) );
  NAND2_X1 U2631 ( .A1(n5761), .A2(n6462), .ZN(n2752) );
  OAI21_X1 U2632 ( .B1(n6086), .B2(n2463), .A(n2753), .ZN(n2750) );
  AOI22_X1 U2633 ( .A1(n5755), .A2(n6398), .B1(n5752), .B2(n6430), .ZN(n2753)
         );
  NAND2_X1 U2634 ( .A1(n2754), .A2(n2755), .ZN(n2749) );
  AOI22_X1 U2635 ( .A1(n5749), .A2(n2820), .B1(n5746), .B2(n6526), .ZN(n2755)
         );
  AOI22_X1 U2636 ( .A1(n5743), .A2(n6366), .B1(n5740), .B2(n6249), .ZN(n2754)
         );
  AOI22_X1 U2638 ( .A1(n5735), .A2(n6566), .B1(n5734), .B2(n6313), .ZN(n2759)
         );
  AOI22_X1 U2639 ( .A1(n5731), .A2(n6150), .B1(n5728), .B2(n6598), .ZN(n2758)
         );
  AOI22_X1 U2640 ( .A1(n5725), .A2(n2235), .B1(n5722), .B2(n2352), .ZN(n2757)
         );
  AOI22_X1 U2641 ( .A1(n5717), .A2(n630), .B1(n5716), .B2(n470), .ZN(n2756) );
  NOR4_X1 U2642 ( .A1(n2760), .A2(n2761), .A3(n2762), .A4(n2763), .ZN(n2746)
         );
  NAND2_X1 U2643 ( .A1(n2764), .A2(n2765), .ZN(n2763) );
  AOI22_X1 U2644 ( .A1(n2491), .A2(n406), .B1(n5709), .B2(n6182), .ZN(n2765)
         );
  AOI22_X1 U2645 ( .A1(n2493), .A2(n6281), .B1(n5458), .B2(OUT1[21]), .ZN(
        n2764) );
  NAND2_X1 U2646 ( .A1(n2766), .A2(n2767), .ZN(n2762) );
  AOI22_X1 U2647 ( .A1(n5704), .A2(n438), .B1(n5701), .B2(n6118), .ZN(n2767)
         );
  AOI22_X1 U2648 ( .A1(n5698), .A2(n6214), .B1(n5695), .B2(n566), .ZN(n2766)
         );
  NAND2_X1 U2649 ( .A1(n2768), .A2(n2769), .ZN(n2761) );
  AOI22_X1 U2650 ( .A1(n5691), .A2(n694), .B1(n5689), .B2(n662), .ZN(n2769) );
  AOI22_X1 U2651 ( .A1(n5686), .A2(n726), .B1(n2505), .B2(n598), .ZN(n2768) );
  NAND2_X1 U2652 ( .A1(n2770), .A2(n2771), .ZN(n2760) );
  AOI22_X1 U2653 ( .A1(n5680), .A2(n502), .B1(n5677), .B2(n374), .ZN(n2771) );
  AOI22_X1 U2654 ( .A1(n5674), .A2(n534), .B1(n5671), .B2(n342), .ZN(n2770) );
  NAND2_X1 U2655 ( .A1(n2772), .A2(n2773), .ZN(n3218) );
  NOR4_X1 U2656 ( .A1(n2774), .A2(n2775), .A3(n2776), .A4(n2777), .ZN(n2773)
         );
  OAI21_X1 U2657 ( .B1(n1434), .B2(n5763), .A(n2778), .ZN(n2777) );
  NAND2_X1 U2658 ( .A1(n5761), .A2(n6463), .ZN(n2778) );
  OAI21_X1 U2659 ( .B1(n6087), .B2(n2463), .A(n2779), .ZN(n2776) );
  AOI22_X1 U2660 ( .A1(n5755), .A2(n6399), .B1(n5752), .B2(n6431), .ZN(n2779)
         );
  NAND2_X1 U2661 ( .A1(n2780), .A2(n2781), .ZN(n2775) );
  AOI22_X1 U2662 ( .A1(n5749), .A2(n2819), .B1(n5746), .B2(n6527), .ZN(n2781)
         );
  AOI22_X1 U2663 ( .A1(n5743), .A2(n6367), .B1(n5740), .B2(n6250), .ZN(n2780)
         );
  AOI22_X1 U2665 ( .A1(n2477), .A2(n6567), .B1(n5734), .B2(n6314), .ZN(n2785)
         );
  AOI22_X1 U2666 ( .A1(n5731), .A2(n6151), .B1(n5728), .B2(n6599), .ZN(n2784)
         );
  AOI22_X1 U2667 ( .A1(n5725), .A2(n2230), .B1(n5722), .B2(n6335), .ZN(n2783)
         );
  AOI22_X1 U2668 ( .A1(n2483), .A2(n629), .B1(n5716), .B2(n469), .ZN(n2782) );
  NOR4_X1 U2669 ( .A1(n2786), .A2(n2787), .A3(n2788), .A4(n2789), .ZN(n2772)
         );
  NAND2_X1 U2670 ( .A1(n2790), .A2(n2791), .ZN(n2789) );
  AOI22_X1 U2671 ( .A1(n5713), .A2(n405), .B1(n5709), .B2(n6183), .ZN(n2791)
         );
  AOI22_X1 U2672 ( .A1(n5707), .A2(n6282), .B1(n5458), .B2(OUT1[20]), .ZN(
        n2790) );
  NAND2_X1 U2673 ( .A1(n2792), .A2(n2793), .ZN(n2788) );
  AOI22_X1 U2674 ( .A1(n5704), .A2(n437), .B1(n5701), .B2(n6119), .ZN(n2793)
         );
  AOI22_X1 U2675 ( .A1(n5698), .A2(n6215), .B1(n5695), .B2(n565), .ZN(n2792)
         );
  NAND2_X1 U2676 ( .A1(n2794), .A2(n2795), .ZN(n2787) );
  AOI22_X1 U2677 ( .A1(n5691), .A2(n693), .B1(n5689), .B2(n661), .ZN(n2795) );
  AOI22_X1 U2678 ( .A1(n5686), .A2(n725), .B1(n2505), .B2(n597), .ZN(n2794) );
  NAND2_X1 U2679 ( .A1(n2796), .A2(n2797), .ZN(n2786) );
  AOI22_X1 U2680 ( .A1(n5680), .A2(n501), .B1(n5677), .B2(n373), .ZN(n2797) );
  AOI22_X1 U2681 ( .A1(n5674), .A2(n533), .B1(n5671), .B2(n341), .ZN(n2796) );
  NAND2_X1 U2682 ( .A1(n2798), .A2(n2799), .ZN(n3217) );
  NOR4_X1 U2683 ( .A1(n2800), .A2(n2801), .A3(n2802), .A4(n2803), .ZN(n2799)
         );
  OAI21_X1 U2684 ( .B1(n1435), .B2(n5763), .A(n2804), .ZN(n2803) );
  NAND2_X1 U2685 ( .A1(n5761), .A2(n6464), .ZN(n2804) );
  OAI21_X1 U2686 ( .B1(n6088), .B2(n2463), .A(n2805), .ZN(n2802) );
  AOI22_X1 U2687 ( .A1(n5755), .A2(n6400), .B1(n5752), .B2(n6432), .ZN(n2805)
         );
  NAND2_X1 U2688 ( .A1(n2806), .A2(n2831), .ZN(n2801) );
  AOI22_X1 U2689 ( .A1(n5749), .A2(n2818), .B1(n5746), .B2(n6528), .ZN(n2831)
         );
  AOI22_X1 U2690 ( .A1(n5743), .A2(n6368), .B1(n5740), .B2(n6251), .ZN(n2806)
         );
  AOI22_X1 U2692 ( .A1(n2477), .A2(n6568), .B1(n5734), .B2(n6315), .ZN(n2835)
         );
  AOI22_X1 U2693 ( .A1(n5731), .A2(n6152), .B1(n5728), .B2(n6600), .ZN(n2834)
         );
  AOI22_X1 U2694 ( .A1(n5725), .A2(n2225), .B1(n5722), .B2(n6336), .ZN(n2833)
         );
  AOI22_X1 U2695 ( .A1(n2483), .A2(n628), .B1(n5716), .B2(n468), .ZN(n2832) );
  NOR4_X1 U2696 ( .A1(n2836), .A2(n2837), .A3(n2838), .A4(n2839), .ZN(n2798)
         );
  NAND2_X1 U2697 ( .A1(n2840), .A2(n2841), .ZN(n2839) );
  AOI22_X1 U2698 ( .A1(n5713), .A2(n404), .B1(n5709), .B2(n6184), .ZN(n2841)
         );
  AOI22_X1 U2699 ( .A1(n5707), .A2(n6283), .B1(n5939), .B2(OUT1[19]), .ZN(
        n2840) );
  NAND2_X1 U2700 ( .A1(n2842), .A2(n2843), .ZN(n2838) );
  AOI22_X1 U2701 ( .A1(n5704), .A2(n436), .B1(n5701), .B2(n6120), .ZN(n2843)
         );
  AOI22_X1 U2702 ( .A1(n5698), .A2(n6216), .B1(n5695), .B2(n564), .ZN(n2842)
         );
  NAND2_X1 U2703 ( .A1(n2844), .A2(n2845), .ZN(n2837) );
  AOI22_X1 U2704 ( .A1(n5691), .A2(n692), .B1(n5689), .B2(n660), .ZN(n2845) );
  AOI22_X1 U2705 ( .A1(n5686), .A2(n724), .B1(n2505), .B2(n596), .ZN(n2844) );
  NAND2_X1 U2706 ( .A1(n2846), .A2(n2847), .ZN(n2836) );
  AOI22_X1 U2707 ( .A1(n5680), .A2(n500), .B1(n5677), .B2(n372), .ZN(n2847) );
  AOI22_X1 U2708 ( .A1(n5674), .A2(n532), .B1(n5671), .B2(n340), .ZN(n2846) );
  NAND2_X1 U2709 ( .A1(n2848), .A2(n2849), .ZN(n3216) );
  NOR4_X1 U2710 ( .A1(n2850), .A2(n2851), .A3(n2852), .A4(n2853), .ZN(n2849)
         );
  OAI21_X1 U2711 ( .B1(n1436), .B2(n5763), .A(n2854), .ZN(n2853) );
  NAND2_X1 U2712 ( .A1(n5761), .A2(n6465), .ZN(n2854) );
  OAI21_X1 U2713 ( .B1(n6089), .B2(n2463), .A(n2855), .ZN(n2852) );
  AOI22_X1 U2714 ( .A1(n5755), .A2(n6401), .B1(n5752), .B2(n6433), .ZN(n2855)
         );
  NAND2_X1 U2715 ( .A1(n2856), .A2(n2857), .ZN(n2851) );
  AOI22_X1 U2716 ( .A1(n5749), .A2(n2817), .B1(n5746), .B2(n6529), .ZN(n2857)
         );
  AOI22_X1 U2717 ( .A1(n5743), .A2(n6369), .B1(n5740), .B2(n6252), .ZN(n2856)
         );
  AOI22_X1 U2719 ( .A1(n2477), .A2(n6569), .B1(n5734), .B2(n6316), .ZN(n2861)
         );
  AOI22_X1 U2720 ( .A1(n5731), .A2(n6153), .B1(n5728), .B2(n6601), .ZN(n2860)
         );
  AOI22_X1 U2721 ( .A1(n5725), .A2(n2220), .B1(n5722), .B2(n6337), .ZN(n2859)
         );
  AOI22_X1 U2722 ( .A1(n2483), .A2(n627), .B1(n5716), .B2(n467), .ZN(n2858) );
  NOR4_X1 U2723 ( .A1(n2862), .A2(n2863), .A3(n2864), .A4(n2865), .ZN(n2848)
         );
  NAND2_X1 U2724 ( .A1(n2866), .A2(n2867), .ZN(n2865) );
  AOI22_X1 U2725 ( .A1(n5713), .A2(n403), .B1(n5709), .B2(n6185), .ZN(n2867)
         );
  AOI22_X1 U2726 ( .A1(n5707), .A2(n6284), .B1(n5939), .B2(OUT1[18]), .ZN(
        n2866) );
  NAND2_X1 U2727 ( .A1(n2868), .A2(n2869), .ZN(n2864) );
  AOI22_X1 U2728 ( .A1(n5704), .A2(n435), .B1(n5701), .B2(n6121), .ZN(n2869)
         );
  AOI22_X1 U2729 ( .A1(n5698), .A2(n6217), .B1(n5695), .B2(n563), .ZN(n2868)
         );
  NAND2_X1 U2730 ( .A1(n2870), .A2(n2871), .ZN(n2863) );
  AOI22_X1 U2731 ( .A1(n5691), .A2(n691), .B1(n5689), .B2(n659), .ZN(n2871) );
  AOI22_X1 U2732 ( .A1(n5686), .A2(n723), .B1(n2505), .B2(n595), .ZN(n2870) );
  NAND2_X1 U2733 ( .A1(n2872), .A2(n2873), .ZN(n2862) );
  AOI22_X1 U2734 ( .A1(n5680), .A2(n499), .B1(n5677), .B2(n371), .ZN(n2873) );
  AOI22_X1 U2735 ( .A1(n5674), .A2(n531), .B1(n5671), .B2(n339), .ZN(n2872) );
  NAND2_X1 U2736 ( .A1(n2874), .A2(n2875), .ZN(n3215) );
  NOR4_X1 U2737 ( .A1(n2876), .A2(n2877), .A3(n2878), .A4(n2879), .ZN(n2875)
         );
  OAI21_X1 U2738 ( .B1(n1437), .B2(n5763), .A(n2880), .ZN(n2879) );
  NAND2_X1 U2739 ( .A1(n5761), .A2(n6466), .ZN(n2880) );
  OAI21_X1 U2740 ( .B1(n6090), .B2(n2463), .A(n2881), .ZN(n2878) );
  AOI22_X1 U2741 ( .A1(n5755), .A2(n6402), .B1(n5752), .B2(n6434), .ZN(n2881)
         );
  NAND2_X1 U2742 ( .A1(n2882), .A2(n2883), .ZN(n2877) );
  AOI22_X1 U2743 ( .A1(n5749), .A2(n2816), .B1(n5746), .B2(n6530), .ZN(n2883)
         );
  AOI22_X1 U2744 ( .A1(n5743), .A2(n6370), .B1(n5740), .B2(n6253), .ZN(n2882)
         );
  AOI22_X1 U2746 ( .A1(n2477), .A2(n6570), .B1(n5734), .B2(n6317), .ZN(n2887)
         );
  AOI22_X1 U2747 ( .A1(n5731), .A2(n6154), .B1(n5728), .B2(n6602), .ZN(n2886)
         );
  AOI22_X1 U2748 ( .A1(n5725), .A2(n2215), .B1(n5722), .B2(n6338), .ZN(n2885)
         );
  AOI22_X1 U2749 ( .A1(n2483), .A2(n626), .B1(n5716), .B2(n466), .ZN(n2884) );
  NOR4_X1 U2750 ( .A1(n2888), .A2(n2889), .A3(n2890), .A4(n2891), .ZN(n2874)
         );
  NAND2_X1 U2751 ( .A1(n2892), .A2(n2893), .ZN(n2891) );
  AOI22_X1 U2752 ( .A1(n5713), .A2(n402), .B1(n5709), .B2(n6186), .ZN(n2893)
         );
  AOI22_X1 U2753 ( .A1(n5707), .A2(n6285), .B1(n5939), .B2(OUT1[17]), .ZN(
        n2892) );
  NAND2_X1 U2754 ( .A1(n2894), .A2(n2895), .ZN(n2890) );
  AOI22_X1 U2755 ( .A1(n5704), .A2(n434), .B1(n5701), .B2(n6122), .ZN(n2895)
         );
  AOI22_X1 U2756 ( .A1(n5698), .A2(n6218), .B1(n5695), .B2(n562), .ZN(n2894)
         );
  NAND2_X1 U2757 ( .A1(n2896), .A2(n2897), .ZN(n2889) );
  AOI22_X1 U2758 ( .A1(n5691), .A2(n690), .B1(n5689), .B2(n658), .ZN(n2897) );
  AOI22_X1 U2759 ( .A1(n5686), .A2(n722), .B1(n2505), .B2(n594), .ZN(n2896) );
  NAND2_X1 U2760 ( .A1(n2898), .A2(n2899), .ZN(n2888) );
  AOI22_X1 U2761 ( .A1(n5680), .A2(n498), .B1(n5677), .B2(n370), .ZN(n2899) );
  AOI22_X1 U2762 ( .A1(n5674), .A2(n530), .B1(n5671), .B2(n338), .ZN(n2898) );
  NAND2_X1 U2763 ( .A1(n2900), .A2(n2901), .ZN(n3214) );
  NOR4_X1 U2764 ( .A1(n2902), .A2(n2903), .A3(n2904), .A4(n2905), .ZN(n2901)
         );
  OAI21_X1 U2765 ( .B1(n1438), .B2(n5763), .A(n2906), .ZN(n2905) );
  NAND2_X1 U2766 ( .A1(n5761), .A2(n6467), .ZN(n2906) );
  OAI21_X1 U2767 ( .B1(n6091), .B2(n2463), .A(n2907), .ZN(n2904) );
  AOI22_X1 U2768 ( .A1(n5755), .A2(n6403), .B1(n5752), .B2(n6435), .ZN(n2907)
         );
  NAND2_X1 U2769 ( .A1(n2908), .A2(n2909), .ZN(n2903) );
  AOI22_X1 U2770 ( .A1(n5749), .A2(n2815), .B1(n5746), .B2(n6531), .ZN(n2909)
         );
  AOI22_X1 U2771 ( .A1(n5743), .A2(n6371), .B1(n5740), .B2(n6254), .ZN(n2908)
         );
  AOI22_X1 U2773 ( .A1(n2477), .A2(n6571), .B1(n5734), .B2(n6318), .ZN(n2913)
         );
  AOI22_X1 U2774 ( .A1(n5731), .A2(n6155), .B1(n5728), .B2(n6603), .ZN(n2912)
         );
  AOI22_X1 U2775 ( .A1(n5725), .A2(n2210), .B1(n5722), .B2(n6339), .ZN(n2911)
         );
  AOI22_X1 U2776 ( .A1(n2483), .A2(n625), .B1(n5716), .B2(n465), .ZN(n2910) );
  NOR4_X1 U2777 ( .A1(n2914), .A2(n2915), .A3(n2916), .A4(n2917), .ZN(n2900)
         );
  NAND2_X1 U2778 ( .A1(n2918), .A2(n2919), .ZN(n2917) );
  AOI22_X1 U2779 ( .A1(n5713), .A2(n401), .B1(n5709), .B2(n6187), .ZN(n2919)
         );
  AOI22_X1 U2780 ( .A1(n5707), .A2(n6286), .B1(n5939), .B2(OUT1[16]), .ZN(
        n2918) );
  NAND2_X1 U2781 ( .A1(n2920), .A2(n2921), .ZN(n2916) );
  AOI22_X1 U2782 ( .A1(n5704), .A2(n433), .B1(n5701), .B2(n6123), .ZN(n2921)
         );
  AOI22_X1 U2783 ( .A1(n5698), .A2(n6219), .B1(n5695), .B2(n561), .ZN(n2920)
         );
  NAND2_X1 U2784 ( .A1(n2922), .A2(n2923), .ZN(n2915) );
  AOI22_X1 U2785 ( .A1(n5691), .A2(n689), .B1(n5689), .B2(n657), .ZN(n2923) );
  AOI22_X1 U2786 ( .A1(n5686), .A2(n721), .B1(n2505), .B2(n593), .ZN(n2922) );
  NAND2_X1 U2787 ( .A1(n2924), .A2(n2925), .ZN(n2914) );
  AOI22_X1 U2788 ( .A1(n5680), .A2(n497), .B1(n5677), .B2(n369), .ZN(n2925) );
  AOI22_X1 U2789 ( .A1(n5674), .A2(n529), .B1(n5671), .B2(n337), .ZN(n2924) );
  NAND2_X1 U2790 ( .A1(n2926), .A2(n2927), .ZN(n3213) );
  NOR4_X1 U2791 ( .A1(n2928), .A2(n2929), .A3(n2930), .A4(n2931), .ZN(n2927)
         );
  OAI21_X1 U2792 ( .B1(n1439), .B2(n5763), .A(n2932), .ZN(n2931) );
  NAND2_X1 U2793 ( .A1(n5761), .A2(n6468), .ZN(n2932) );
  OAI21_X1 U2794 ( .B1(n5507), .B2(n2463), .A(n2933), .ZN(n2930) );
  AOI22_X1 U2795 ( .A1(n5755), .A2(n6404), .B1(n5752), .B2(n6436), .ZN(n2933)
         );
  NAND2_X1 U2796 ( .A1(n2934), .A2(n2935), .ZN(n2929) );
  AOI22_X1 U2797 ( .A1(n5749), .A2(n2814), .B1(n5746), .B2(n6532), .ZN(n2935)
         );
  AOI22_X1 U2798 ( .A1(n5743), .A2(n6372), .B1(n5740), .B2(n6255), .ZN(n2934)
         );
  AOI22_X1 U2800 ( .A1(n2477), .A2(n6572), .B1(n5734), .B2(n6319), .ZN(n2939)
         );
  AOI22_X1 U2801 ( .A1(n5731), .A2(n6156), .B1(n5728), .B2(n6604), .ZN(n2938)
         );
  AOI22_X1 U2802 ( .A1(n5725), .A2(n2205), .B1(n5722), .B2(n6340), .ZN(n2937)
         );
  AOI22_X1 U2803 ( .A1(n2483), .A2(n624), .B1(n5716), .B2(n464), .ZN(n2936) );
  NOR4_X1 U2804 ( .A1(n2940), .A2(n2941), .A3(n2942), .A4(n2943), .ZN(n2926)
         );
  NAND2_X1 U2805 ( .A1(n2944), .A2(n2945), .ZN(n2943) );
  AOI22_X1 U2806 ( .A1(n5713), .A2(n400), .B1(n5709), .B2(n6188), .ZN(n2945)
         );
  AOI22_X1 U2807 ( .A1(n5707), .A2(n6287), .B1(n5939), .B2(OUT1[15]), .ZN(
        n2944) );
  NAND2_X1 U2808 ( .A1(n2946), .A2(n2947), .ZN(n2942) );
  AOI22_X1 U2809 ( .A1(n5704), .A2(n432), .B1(n5701), .B2(n6124), .ZN(n2947)
         );
  AOI22_X1 U2810 ( .A1(n5698), .A2(n6220), .B1(n5695), .B2(n560), .ZN(n2946)
         );
  NAND2_X1 U2811 ( .A1(n2948), .A2(n2949), .ZN(n2941) );
  AOI22_X1 U2812 ( .A1(n5691), .A2(n688), .B1(n5689), .B2(n656), .ZN(n2949) );
  AOI22_X1 U2813 ( .A1(n5686), .A2(n720), .B1(n2505), .B2(n592), .ZN(n2948) );
  NAND2_X1 U2814 ( .A1(n2950), .A2(n2951), .ZN(n2940) );
  AOI22_X1 U2815 ( .A1(n5680), .A2(n496), .B1(n5677), .B2(n368), .ZN(n2951) );
  AOI22_X1 U2816 ( .A1(n5674), .A2(n528), .B1(n5671), .B2(n336), .ZN(n2950) );
  NAND2_X1 U2817 ( .A1(n2952), .A2(n2953), .ZN(n3212) );
  NOR4_X1 U2818 ( .A1(n2954), .A2(n2955), .A3(n2956), .A4(n2957), .ZN(n2953)
         );
  OAI21_X1 U2819 ( .B1(n1440), .B2(n5763), .A(n2958), .ZN(n2957) );
  NAND2_X1 U2820 ( .A1(n5761), .A2(n6469), .ZN(n2958) );
  OAI21_X1 U2821 ( .B1(n6093), .B2(n2463), .A(n2959), .ZN(n2956) );
  AOI22_X1 U2822 ( .A1(n5755), .A2(n6405), .B1(n5752), .B2(n6437), .ZN(n2959)
         );
  NAND2_X1 U2823 ( .A1(n2960), .A2(n2961), .ZN(n2955) );
  AOI22_X1 U2824 ( .A1(n5749), .A2(n2813), .B1(n5746), .B2(n6533), .ZN(n2961)
         );
  AOI22_X1 U2825 ( .A1(n5743), .A2(n6373), .B1(n5740), .B2(n6256), .ZN(n2960)
         );
  AOI22_X1 U2827 ( .A1(n2477), .A2(n6573), .B1(n5734), .B2(n6320), .ZN(n2965)
         );
  AOI22_X1 U2828 ( .A1(n5731), .A2(n6157), .B1(n5728), .B2(n6605), .ZN(n2964)
         );
  AOI22_X1 U2829 ( .A1(n5725), .A2(n2200), .B1(n5722), .B2(n6341), .ZN(n2963)
         );
  AOI22_X1 U2830 ( .A1(n2483), .A2(n623), .B1(n5716), .B2(n463), .ZN(n2962) );
  NOR4_X1 U2831 ( .A1(n2966), .A2(n2967), .A3(n2968), .A4(n2969), .ZN(n2952)
         );
  NAND2_X1 U2832 ( .A1(n2970), .A2(n2971), .ZN(n2969) );
  AOI22_X1 U2833 ( .A1(n5713), .A2(n399), .B1(n5709), .B2(n6189), .ZN(n2971)
         );
  AOI22_X1 U2834 ( .A1(n5707), .A2(n6288), .B1(n5939), .B2(OUT1[14]), .ZN(
        n2970) );
  NAND2_X1 U2835 ( .A1(n2972), .A2(n2973), .ZN(n2968) );
  AOI22_X1 U2836 ( .A1(n5704), .A2(n431), .B1(n5701), .B2(n6125), .ZN(n2973)
         );
  AOI22_X1 U2837 ( .A1(n5698), .A2(n6221), .B1(n5695), .B2(n559), .ZN(n2972)
         );
  NAND2_X1 U2838 ( .A1(n2974), .A2(n2975), .ZN(n2967) );
  AOI22_X1 U2839 ( .A1(n5691), .A2(n687), .B1(n5689), .B2(n655), .ZN(n2975) );
  AOI22_X1 U2840 ( .A1(n5686), .A2(n719), .B1(n2505), .B2(n591), .ZN(n2974) );
  NAND2_X1 U2841 ( .A1(n2976), .A2(n2977), .ZN(n2966) );
  AOI22_X1 U2842 ( .A1(n5680), .A2(n495), .B1(n5677), .B2(n367), .ZN(n2977) );
  AOI22_X1 U2843 ( .A1(n5674), .A2(n527), .B1(n5671), .B2(n335), .ZN(n2976) );
  NAND2_X1 U2844 ( .A1(n2978), .A2(n2979), .ZN(n3211) );
  NOR4_X1 U2845 ( .A1(n2980), .A2(n2981), .A3(n2982), .A4(n2983), .ZN(n2979)
         );
  OAI21_X1 U2846 ( .B1(n1441), .B2(n5763), .A(n2984), .ZN(n2983) );
  NAND2_X1 U2847 ( .A1(n5761), .A2(n6470), .ZN(n2984) );
  OAI21_X1 U2848 ( .B1(n6094), .B2(n2463), .A(n2985), .ZN(n2982) );
  AOI22_X1 U2849 ( .A1(n5755), .A2(n6406), .B1(n5752), .B2(n6438), .ZN(n2985)
         );
  NAND2_X1 U2850 ( .A1(n2986), .A2(n2987), .ZN(n2981) );
  AOI22_X1 U2851 ( .A1(n5749), .A2(n2812), .B1(n5746), .B2(n6534), .ZN(n2987)
         );
  AOI22_X1 U2852 ( .A1(n5743), .A2(n6374), .B1(n5740), .B2(n6257), .ZN(n2986)
         );
  AOI22_X1 U2854 ( .A1(n2477), .A2(n6574), .B1(n5734), .B2(n6321), .ZN(n2991)
         );
  AOI22_X1 U2855 ( .A1(n5731), .A2(n6158), .B1(n5728), .B2(n6606), .ZN(n2990)
         );
  AOI22_X1 U2856 ( .A1(n5725), .A2(n2195), .B1(n5722), .B2(n6342), .ZN(n2989)
         );
  AOI22_X1 U2857 ( .A1(n2483), .A2(n622), .B1(n5716), .B2(n462), .ZN(n2988) );
  NOR4_X1 U2858 ( .A1(n2992), .A2(n2993), .A3(n2994), .A4(n2995), .ZN(n2978)
         );
  NAND2_X1 U2859 ( .A1(n2996), .A2(n2997), .ZN(n2995) );
  AOI22_X1 U2860 ( .A1(n5713), .A2(n398), .B1(n5709), .B2(n6190), .ZN(n2997)
         );
  AOI22_X1 U2861 ( .A1(n5707), .A2(n6289), .B1(n5939), .B2(OUT1[13]), .ZN(
        n2996) );
  NAND2_X1 U2862 ( .A1(n2998), .A2(n2999), .ZN(n2994) );
  AOI22_X1 U2863 ( .A1(n2496), .A2(n430), .B1(n5701), .B2(n6126), .ZN(n2999)
         );
  AOI22_X1 U2864 ( .A1(n5698), .A2(n6222), .B1(n5695), .B2(n558), .ZN(n2998)
         );
  NAND2_X1 U2865 ( .A1(n3000), .A2(n3001), .ZN(n2993) );
  AOI22_X1 U2866 ( .A1(n5691), .A2(n686), .B1(n5689), .B2(n654), .ZN(n3001) );
  AOI22_X1 U2867 ( .A1(n5686), .A2(n718), .B1(n2505), .B2(n590), .ZN(n3000) );
  NAND2_X1 U2868 ( .A1(n3002), .A2(n3003), .ZN(n2992) );
  AOI22_X1 U2869 ( .A1(n2508), .A2(n494), .B1(n5677), .B2(n366), .ZN(n3003) );
  AOI22_X1 U2870 ( .A1(n5674), .A2(n526), .B1(n5671), .B2(n334), .ZN(n3002) );
  NAND2_X1 U2871 ( .A1(n3004), .A2(n3005), .ZN(n3210) );
  NOR4_X1 U2872 ( .A1(n3006), .A2(n3007), .A3(n3008), .A4(n3009), .ZN(n3005)
         );
  OAI21_X1 U2873 ( .B1(n1442), .B2(n5763), .A(n3010), .ZN(n3009) );
  NAND2_X1 U2874 ( .A1(n5761), .A2(n6471), .ZN(n3010) );
  OAI21_X1 U2875 ( .B1(n6095), .B2(n2463), .A(n3011), .ZN(n3008) );
  AOI22_X1 U2876 ( .A1(n2465), .A2(n6407), .B1(n5752), .B2(n6439), .ZN(n3011)
         );
  NAND2_X1 U2877 ( .A1(n3012), .A2(n3013), .ZN(n3007) );
  AOI22_X1 U2878 ( .A1(n2469), .A2(n2811), .B1(n5746), .B2(n6535), .ZN(n3013)
         );
  AOI22_X1 U2879 ( .A1(n2471), .A2(n6375), .B1(n5740), .B2(n6258), .ZN(n3012)
         );
  AOI22_X1 U2881 ( .A1(n2477), .A2(n6575), .B1(n5734), .B2(n6322), .ZN(n3017)
         );
  AOI22_X1 U2882 ( .A1(n2479), .A2(n6159), .B1(n5728), .B2(n6607), .ZN(n3016)
         );
  AOI22_X1 U2883 ( .A1(n2481), .A2(n2190), .B1(n5722), .B2(n6343), .ZN(n3015)
         );
  AOI22_X1 U2884 ( .A1(n2483), .A2(n621), .B1(n5716), .B2(n461), .ZN(n3014) );
  NOR4_X1 U2885 ( .A1(n3018), .A2(n3019), .A3(n3020), .A4(n3021), .ZN(n3004)
         );
  NAND2_X1 U2886 ( .A1(n3022), .A2(n3023), .ZN(n3021) );
  AOI22_X1 U2887 ( .A1(n5713), .A2(n397), .B1(n5709), .B2(n6191), .ZN(n3023)
         );
  AOI22_X1 U2888 ( .A1(n5707), .A2(n6290), .B1(n5939), .B2(OUT1[12]), .ZN(
        n3022) );
  NAND2_X1 U2889 ( .A1(n3024), .A2(n3025), .ZN(n3020) );
  AOI22_X1 U2890 ( .A1(n5704), .A2(n429), .B1(n5701), .B2(n6127), .ZN(n3025)
         );
  AOI22_X1 U2891 ( .A1(n2498), .A2(n6223), .B1(n5695), .B2(n557), .ZN(n3024)
         );
  NAND2_X1 U2892 ( .A1(n3026), .A2(n3027), .ZN(n3019) );
  AOI22_X1 U2893 ( .A1(n5691), .A2(n685), .B1(n5689), .B2(n653), .ZN(n3027) );
  AOI22_X1 U2894 ( .A1(n2504), .A2(n717), .B1(n2505), .B2(n589), .ZN(n3026) );
  NAND2_X1 U2895 ( .A1(n3028), .A2(n3029), .ZN(n3018) );
  AOI22_X1 U2896 ( .A1(n5680), .A2(n493), .B1(n5677), .B2(n365), .ZN(n3029) );
  AOI22_X1 U2897 ( .A1(n2510), .A2(n525), .B1(n5671), .B2(n333), .ZN(n3028) );
  NAND2_X1 U2898 ( .A1(n3030), .A2(n3031), .ZN(n3209) );
  NOR4_X1 U2899 ( .A1(n3032), .A2(n3033), .A3(n3034), .A4(n3035), .ZN(n3031)
         );
  OAI21_X1 U2900 ( .B1(n1443), .B2(n5763), .A(n3036), .ZN(n3035) );
  NAND2_X1 U2901 ( .A1(n5761), .A2(n6472), .ZN(n3036) );
  OAI21_X1 U2902 ( .B1(n6096), .B2(n2463), .A(n3037), .ZN(n3034) );
  AOI22_X1 U2903 ( .A1(n5755), .A2(n6408), .B1(n5752), .B2(n6440), .ZN(n3037)
         );
  NAND2_X1 U2904 ( .A1(n3038), .A2(n3039), .ZN(n3033) );
  AOI22_X1 U2905 ( .A1(n5749), .A2(n2810), .B1(n5746), .B2(n6536), .ZN(n3039)
         );
  AOI22_X1 U2906 ( .A1(n5743), .A2(n6376), .B1(n5740), .B2(n6259), .ZN(n3038)
         );
  AOI22_X1 U2908 ( .A1(n5735), .A2(n6576), .B1(n5734), .B2(n6323), .ZN(n3043)
         );
  AOI22_X1 U2909 ( .A1(n5731), .A2(n6160), .B1(n5728), .B2(n6608), .ZN(n3042)
         );
  AOI22_X1 U2910 ( .A1(n5725), .A2(n2185), .B1(n5722), .B2(n6344), .ZN(n3041)
         );
  AOI22_X1 U2911 ( .A1(n5717), .A2(n620), .B1(n5716), .B2(n460), .ZN(n3040) );
  NOR4_X1 U2912 ( .A1(n3044), .A2(n3045), .A3(n3046), .A4(n3047), .ZN(n3030)
         );
  NAND2_X1 U2913 ( .A1(n3048), .A2(n3049), .ZN(n3047) );
  AOI22_X1 U2914 ( .A1(n5713), .A2(n396), .B1(n5709), .B2(n6192), .ZN(n3049)
         );
  AOI22_X1 U2915 ( .A1(n5707), .A2(n6291), .B1(n5939), .B2(OUT1[11]), .ZN(
        n3048) );
  NAND2_X1 U2916 ( .A1(n3050), .A2(n3051), .ZN(n3046) );
  AOI22_X1 U2917 ( .A1(n5704), .A2(n428), .B1(n5701), .B2(n6128), .ZN(n3051)
         );
  AOI22_X1 U2918 ( .A1(n5698), .A2(n6224), .B1(n5695), .B2(n556), .ZN(n3050)
         );
  NAND2_X1 U2919 ( .A1(n3052), .A2(n3053), .ZN(n3045) );
  AOI22_X1 U2920 ( .A1(n5691), .A2(n684), .B1(n5689), .B2(n652), .ZN(n3053) );
  AOI22_X1 U2921 ( .A1(n5686), .A2(n716), .B1(n5681), .B2(n588), .ZN(n3052) );
  NAND2_X1 U2922 ( .A1(n3054), .A2(n3919), .ZN(n3044) );
  AOI22_X1 U2923 ( .A1(n5680), .A2(n492), .B1(n5677), .B2(n364), .ZN(n3919) );
  AOI22_X1 U2924 ( .A1(n5674), .A2(n524), .B1(n5671), .B2(n332), .ZN(n3054) );
  NAND2_X1 U2925 ( .A1(n3920), .A2(n3921), .ZN(n3208) );
  NOR4_X1 U2926 ( .A1(n3922), .A2(n3923), .A3(n3924), .A4(n3925), .ZN(n3921)
         );
  OAI21_X1 U2927 ( .B1(n1444), .B2(n2460), .A(n3926), .ZN(n3925) );
  NAND2_X1 U2928 ( .A1(n2462), .A2(n6473), .ZN(n3926) );
  OAI21_X1 U2929 ( .B1(n6097), .B2(n2463), .A(n3927), .ZN(n3924) );
  AOI22_X1 U2930 ( .A1(n5755), .A2(n6409), .B1(n2466), .B2(n6441), .ZN(n3927)
         );
  NAND2_X1 U2931 ( .A1(n3928), .A2(n3929), .ZN(n3923) );
  AOI22_X1 U2932 ( .A1(n5749), .A2(n2809), .B1(n2470), .B2(n6537), .ZN(n3929)
         );
  AOI22_X1 U2933 ( .A1(n5743), .A2(n6377), .B1(n2472), .B2(n6260), .ZN(n3928)
         );
  AOI22_X1 U2935 ( .A1(n5735), .A2(n6577), .B1(n2478), .B2(n6324), .ZN(n3933)
         );
  AOI22_X1 U2936 ( .A1(n5731), .A2(n6161), .B1(n2480), .B2(n6609), .ZN(n3932)
         );
  AOI22_X1 U2937 ( .A1(n5725), .A2(n2180), .B1(n2482), .B2(n6345), .ZN(n3931)
         );
  AOI22_X1 U2938 ( .A1(n5717), .A2(n619), .B1(n2484), .B2(n459), .ZN(n3930) );
  NOR4_X1 U2939 ( .A1(n3934), .A2(n3935), .A3(n3936), .A4(n3937), .ZN(n3920)
         );
  NAND2_X1 U2940 ( .A1(n3938), .A2(n3939), .ZN(n3937) );
  AOI22_X1 U2941 ( .A1(n5713), .A2(n395), .B1(n5709), .B2(n6193), .ZN(n3939)
         );
  AOI22_X1 U2942 ( .A1(n2493), .A2(n6292), .B1(n5939), .B2(OUT1[10]), .ZN(
        n3938) );
  NAND2_X1 U2943 ( .A1(n3940), .A2(n3941), .ZN(n3936) );
  AOI22_X1 U2944 ( .A1(n2496), .A2(n427), .B1(n2497), .B2(n6129), .ZN(n3941)
         );
  AOI22_X1 U2945 ( .A1(n5698), .A2(n6225), .B1(n2499), .B2(n555), .ZN(n3940)
         );
  NAND2_X1 U2946 ( .A1(n3942), .A2(n3943), .ZN(n3935) );
  AOI22_X1 U2947 ( .A1(n5691), .A2(n683), .B1(n2503), .B2(n651), .ZN(n3943) );
  AOI22_X1 U2948 ( .A1(n5686), .A2(n715), .B1(n5681), .B2(n587), .ZN(n3942) );
  NAND2_X1 U2949 ( .A1(n3944), .A2(n3945), .ZN(n3934) );
  AOI22_X1 U2950 ( .A1(n2508), .A2(n491), .B1(n2509), .B2(n363), .ZN(n3945) );
  AOI22_X1 U2951 ( .A1(n5674), .A2(n523), .B1(n2511), .B2(n331), .ZN(n3944) );
  NAND2_X1 U2952 ( .A1(n3946), .A2(n3947), .ZN(n3207) );
  NOR4_X1 U2953 ( .A1(n3948), .A2(n3949), .A3(n3950), .A4(n3951), .ZN(n3947)
         );
  OAI21_X1 U2954 ( .B1(n1445), .B2(n2460), .A(n3952), .ZN(n3951) );
  NAND2_X1 U2955 ( .A1(n2462), .A2(n6474), .ZN(n3952) );
  OAI21_X1 U2956 ( .B1(n5525), .B2(n2463), .A(n3953), .ZN(n3950) );
  AOI22_X1 U2957 ( .A1(n2465), .A2(n6410), .B1(n2466), .B2(n6442), .ZN(n3953)
         );
  NAND2_X1 U2958 ( .A1(n3954), .A2(n3955), .ZN(n3949) );
  AOI22_X1 U2959 ( .A1(n2469), .A2(n2808), .B1(n2470), .B2(n6538), .ZN(n3955)
         );
  AOI22_X1 U2960 ( .A1(n2471), .A2(n6378), .B1(n2472), .B2(n6261), .ZN(n3954)
         );
  AOI22_X1 U2962 ( .A1(n5735), .A2(n6578), .B1(n2478), .B2(n6325), .ZN(n3959)
         );
  AOI22_X1 U2963 ( .A1(n2479), .A2(n6162), .B1(n2480), .B2(n6610), .ZN(n3958)
         );
  AOI22_X1 U2964 ( .A1(n2481), .A2(n2175), .B1(n2482), .B2(n6346), .ZN(n3957)
         );
  AOI22_X1 U2965 ( .A1(n5717), .A2(n618), .B1(n2484), .B2(n458), .ZN(n3956) );
  NOR4_X1 U2966 ( .A1(n3960), .A2(n3961), .A3(n3962), .A4(n3963), .ZN(n3946)
         );
  NAND2_X1 U2967 ( .A1(n3964), .A2(n3965), .ZN(n3963) );
  AOI22_X1 U2968 ( .A1(n2491), .A2(n394), .B1(n5709), .B2(n6194), .ZN(n3965)
         );
  AOI22_X1 U2969 ( .A1(n2493), .A2(n6293), .B1(n5939), .B2(OUT1[9]), .ZN(n3964) );
  NAND2_X1 U2970 ( .A1(n3966), .A2(n3967), .ZN(n3962) );
  AOI22_X1 U2971 ( .A1(n5704), .A2(n426), .B1(n2497), .B2(n6130), .ZN(n3967)
         );
  AOI22_X1 U2972 ( .A1(n2498), .A2(n6226), .B1(n2499), .B2(n554), .ZN(n3966)
         );
  NAND2_X1 U2973 ( .A1(n3968), .A2(n3969), .ZN(n3961) );
  AOI22_X1 U2974 ( .A1(n5691), .A2(n682), .B1(n2503), .B2(n650), .ZN(n3969) );
  AOI22_X1 U2975 ( .A1(n2504), .A2(n714), .B1(n5681), .B2(n586), .ZN(n3968) );
  NAND2_X1 U2976 ( .A1(n3970), .A2(n3971), .ZN(n3960) );
  AOI22_X1 U2977 ( .A1(n5680), .A2(n490), .B1(n2509), .B2(n362), .ZN(n3971) );
  AOI22_X1 U2978 ( .A1(n2510), .A2(n522), .B1(n2511), .B2(n330), .ZN(n3970) );
  NAND2_X1 U2979 ( .A1(n3972), .A2(n3973), .ZN(n3206) );
  NOR4_X1 U2980 ( .A1(n3974), .A2(n3975), .A3(n3976), .A4(n3977), .ZN(n3973)
         );
  OAI21_X1 U2981 ( .B1(n1446), .B2(n2460), .A(n3978), .ZN(n3977) );
  NAND2_X1 U2982 ( .A1(n2462), .A2(n6475), .ZN(n3978) );
  OAI21_X1 U2983 ( .B1(n6099), .B2(n2463), .A(n3979), .ZN(n3976) );
  AOI22_X1 U2984 ( .A1(n2465), .A2(n6411), .B1(n2466), .B2(n6443), .ZN(n3979)
         );
  NAND2_X1 U2985 ( .A1(n3980), .A2(n3981), .ZN(n3975) );
  AOI22_X1 U2986 ( .A1(n2469), .A2(n2807), .B1(n2470), .B2(n6539), .ZN(n3981)
         );
  AOI22_X1 U2987 ( .A1(n2471), .A2(n6379), .B1(n2472), .B2(n6262), .ZN(n3980)
         );
  AOI22_X1 U2989 ( .A1(n5735), .A2(n6579), .B1(n2478), .B2(n6326), .ZN(n3985)
         );
  AOI22_X1 U2990 ( .A1(n2479), .A2(n6163), .B1(n2480), .B2(n6611), .ZN(n3984)
         );
  AOI22_X1 U2991 ( .A1(n2481), .A2(n2170), .B1(n2482), .B2(n6347), .ZN(n3983)
         );
  AOI22_X1 U2992 ( .A1(n5717), .A2(n617), .B1(n2484), .B2(n457), .ZN(n3982) );
  NOR4_X1 U2993 ( .A1(n3986), .A2(n3987), .A3(n3988), .A4(n3989), .ZN(n3972)
         );
  NAND2_X1 U2994 ( .A1(n3990), .A2(n3991), .ZN(n3989) );
  AOI22_X1 U2995 ( .A1(n2491), .A2(n393), .B1(n5709), .B2(n6195), .ZN(n3991)
         );
  AOI22_X1 U2996 ( .A1(n2493), .A2(n6294), .B1(n5939), .B2(OUT1[8]), .ZN(n3990) );
  NAND2_X1 U2997 ( .A1(n3992), .A2(n3993), .ZN(n3988) );
  AOI22_X1 U2998 ( .A1(n2496), .A2(n425), .B1(n2497), .B2(n6131), .ZN(n3993)
         );
  AOI22_X1 U2999 ( .A1(n2498), .A2(n6227), .B1(n2499), .B2(n553), .ZN(n3992)
         );
  NAND2_X1 U3000 ( .A1(n3994), .A2(n3995), .ZN(n3987) );
  AOI22_X1 U3001 ( .A1(n5691), .A2(n681), .B1(n2503), .B2(n649), .ZN(n3995) );
  AOI22_X1 U3002 ( .A1(n2504), .A2(n713), .B1(n5681), .B2(n585), .ZN(n3994) );
  NAND2_X1 U3003 ( .A1(n3996), .A2(n3997), .ZN(n3986) );
  AOI22_X1 U3004 ( .A1(n2508), .A2(n489), .B1(n2509), .B2(n361), .ZN(n3997) );
  AOI22_X1 U3005 ( .A1(n2510), .A2(n521), .B1(n2511), .B2(n329), .ZN(n3996) );
  NAND2_X1 U3006 ( .A1(n4190), .A2(n4191), .ZN(n3205) );
  NOR4_X1 U3007 ( .A1(n4192), .A2(n4193), .A3(n4194), .A4(n4195), .ZN(n4191)
         );
  OAI21_X1 U3008 ( .B1(n1447), .B2(n2460), .A(n4196), .ZN(n4195) );
  NAND2_X1 U3009 ( .A1(n2462), .A2(n6476), .ZN(n4196) );
  OAI21_X1 U3010 ( .B1(n6100), .B2(n2463), .A(n4197), .ZN(n4194) );
  AOI22_X1 U3011 ( .A1(n2465), .A2(n6412), .B1(n2466), .B2(n6444), .ZN(n4197)
         );
  NAND2_X1 U3012 ( .A1(n4198), .A2(n4199), .ZN(n4193) );
  AOI22_X1 U3013 ( .A1(n2469), .A2(n6548), .B1(n2470), .B2(n6540), .ZN(n4199)
         );
  AOI22_X1 U3014 ( .A1(n2471), .A2(n6380), .B1(n2472), .B2(n6263), .ZN(n4198)
         );
  AOI22_X1 U3016 ( .A1(n5735), .A2(n6580), .B1(n2478), .B2(n6327), .ZN(n4203)
         );
  AOI22_X1 U3017 ( .A1(n2479), .A2(n6164), .B1(n2480), .B2(n6612), .ZN(n4202)
         );
  AOI22_X1 U3018 ( .A1(n2481), .A2(n2165), .B1(n2482), .B2(n6348), .ZN(n4201)
         );
  AOI22_X1 U3019 ( .A1(n5717), .A2(n616), .B1(n2484), .B2(n456), .ZN(n4200) );
  NOR4_X1 U3020 ( .A1(n4204), .A2(n4205), .A3(n4206), .A4(n4207), .ZN(n4190)
         );
  NAND2_X1 U3021 ( .A1(n4208), .A2(n4209), .ZN(n4207) );
  AOI22_X1 U3022 ( .A1(n2491), .A2(n392), .B1(n5709), .B2(n6196), .ZN(n4209)
         );
  AOI22_X1 U3023 ( .A1(n2493), .A2(n6295), .B1(n5939), .B2(OUT1[7]), .ZN(n4208) );
  NAND2_X1 U3024 ( .A1(n4210), .A2(n4211), .ZN(n4206) );
  AOI22_X1 U3025 ( .A1(n2496), .A2(n424), .B1(n2497), .B2(n6132), .ZN(n4211)
         );
  AOI22_X1 U3026 ( .A1(n2498), .A2(n6228), .B1(n2499), .B2(n552), .ZN(n4210)
         );
  NAND2_X1 U3027 ( .A1(n4212), .A2(n4213), .ZN(n4205) );
  AOI22_X1 U3028 ( .A1(n5691), .A2(n680), .B1(n2503), .B2(n648), .ZN(n4213) );
  AOI22_X1 U3029 ( .A1(n2504), .A2(n712), .B1(n5681), .B2(n584), .ZN(n4212) );
  NAND2_X1 U3030 ( .A1(n4214), .A2(n4215), .ZN(n4204) );
  AOI22_X1 U3031 ( .A1(n2508), .A2(n488), .B1(n2509), .B2(n360), .ZN(n4215) );
  AOI22_X1 U3032 ( .A1(n2510), .A2(n520), .B1(n2511), .B2(n328), .ZN(n4214) );
  NAND2_X1 U3033 ( .A1(n4216), .A2(n4217), .ZN(n3204) );
  NOR4_X1 U3034 ( .A1(n4218), .A2(n4219), .A3(n4220), .A4(n4221), .ZN(n4217)
         );
  OAI21_X1 U3035 ( .B1(n1448), .B2(n2460), .A(n4222), .ZN(n4221) );
  NAND2_X1 U3036 ( .A1(n2462), .A2(n6477), .ZN(n4222) );
  OAI21_X1 U3037 ( .B1(n6101), .B2(n2463), .A(n4223), .ZN(n4220) );
  AOI22_X1 U3038 ( .A1(n2465), .A2(n6413), .B1(n2466), .B2(n6445), .ZN(n4223)
         );
  NAND2_X1 U3039 ( .A1(n4224), .A2(n4225), .ZN(n4219) );
  AOI22_X1 U3040 ( .A1(n2469), .A2(n6549), .B1(n2470), .B2(n6541), .ZN(n4225)
         );
  AOI22_X1 U3041 ( .A1(n2471), .A2(n6381), .B1(n2472), .B2(n6264), .ZN(n4224)
         );
  AOI22_X1 U3043 ( .A1(n5735), .A2(n6581), .B1(n2478), .B2(n6328), .ZN(n4229)
         );
  AOI22_X1 U3044 ( .A1(n2479), .A2(n6165), .B1(n2480), .B2(n6613), .ZN(n4228)
         );
  AOI22_X1 U3045 ( .A1(n2481), .A2(n2160), .B1(n2482), .B2(n6349), .ZN(n4227)
         );
  AOI22_X1 U3046 ( .A1(n5717), .A2(n615), .B1(n2484), .B2(n455), .ZN(n4226) );
  NOR4_X1 U3047 ( .A1(n4230), .A2(n4231), .A3(n4232), .A4(n4233), .ZN(n4216)
         );
  NAND2_X1 U3048 ( .A1(n4234), .A2(n4235), .ZN(n4233) );
  AOI22_X1 U3049 ( .A1(n2491), .A2(n391), .B1(n5709), .B2(n6197), .ZN(n4235)
         );
  AOI22_X1 U3050 ( .A1(n2493), .A2(n6296), .B1(n5939), .B2(OUT1[6]), .ZN(n4234) );
  NAND2_X1 U3051 ( .A1(n4236), .A2(n4237), .ZN(n4232) );
  AOI22_X1 U3052 ( .A1(n2496), .A2(n423), .B1(n2497), .B2(n6133), .ZN(n4237)
         );
  AOI22_X1 U3053 ( .A1(n2498), .A2(n6229), .B1(n2499), .B2(n551), .ZN(n4236)
         );
  NAND2_X1 U3054 ( .A1(n4238), .A2(n4239), .ZN(n4231) );
  AOI22_X1 U3055 ( .A1(n5691), .A2(n679), .B1(n2503), .B2(n647), .ZN(n4239) );
  AOI22_X1 U3056 ( .A1(n2504), .A2(n711), .B1(n5681), .B2(n583), .ZN(n4238) );
  NAND2_X1 U3057 ( .A1(n4240), .A2(n4241), .ZN(n4230) );
  AOI22_X1 U3058 ( .A1(n2508), .A2(n487), .B1(n2509), .B2(n359), .ZN(n4241) );
  AOI22_X1 U3059 ( .A1(n2510), .A2(n519), .B1(n2511), .B2(n327), .ZN(n4240) );
  NAND2_X1 U3060 ( .A1(n4242), .A2(n4243), .ZN(n3203) );
  NOR4_X1 U3061 ( .A1(n4244), .A2(n4245), .A3(n4246), .A4(n4247), .ZN(n4243)
         );
  OAI21_X1 U3062 ( .B1(n1449), .B2(n2460), .A(n4248), .ZN(n4247) );
  NAND2_X1 U3063 ( .A1(n2462), .A2(n6478), .ZN(n4248) );
  OAI21_X1 U3064 ( .B1(n6102), .B2(n2463), .A(n4249), .ZN(n4246) );
  AOI22_X1 U3065 ( .A1(n2465), .A2(n6414), .B1(n2466), .B2(n6446), .ZN(n4249)
         );
  NAND2_X1 U3066 ( .A1(n4250), .A2(n4251), .ZN(n4245) );
  AOI22_X1 U3067 ( .A1(n2469), .A2(n6550), .B1(n2470), .B2(n6542), .ZN(n4251)
         );
  AOI22_X1 U3068 ( .A1(n2471), .A2(n6382), .B1(n2472), .B2(n6265), .ZN(n4250)
         );
  AOI22_X1 U3070 ( .A1(n5735), .A2(n6582), .B1(n2478), .B2(n6329), .ZN(n4255)
         );
  AOI22_X1 U3071 ( .A1(n2479), .A2(n6166), .B1(n2480), .B2(n6614), .ZN(n4254)
         );
  AOI22_X1 U3072 ( .A1(n2481), .A2(n2155), .B1(n2482), .B2(n6350), .ZN(n4253)
         );
  AOI22_X1 U3073 ( .A1(n5717), .A2(n614), .B1(n2484), .B2(n454), .ZN(n4252) );
  NOR4_X1 U3074 ( .A1(n4256), .A2(n4257), .A3(n4258), .A4(n4259), .ZN(n4242)
         );
  NAND2_X1 U3075 ( .A1(n4260), .A2(n4261), .ZN(n4259) );
  AOI22_X1 U3076 ( .A1(n2491), .A2(n390), .B1(n5709), .B2(n6198), .ZN(n4261)
         );
  AOI22_X1 U3077 ( .A1(n2493), .A2(n6297), .B1(n5939), .B2(OUT1[5]), .ZN(n4260) );
  NAND2_X1 U3078 ( .A1(n4262), .A2(n4263), .ZN(n4258) );
  AOI22_X1 U3079 ( .A1(n2496), .A2(n422), .B1(n2497), .B2(n6134), .ZN(n4263)
         );
  AOI22_X1 U3080 ( .A1(n2498), .A2(n6230), .B1(n2499), .B2(n550), .ZN(n4262)
         );
  NAND2_X1 U3081 ( .A1(n4264), .A2(n4265), .ZN(n4257) );
  AOI22_X1 U3082 ( .A1(n5691), .A2(n678), .B1(n2503), .B2(n646), .ZN(n4265) );
  AOI22_X1 U3083 ( .A1(n2504), .A2(n710), .B1(n5681), .B2(n582), .ZN(n4264) );
  NAND2_X1 U3084 ( .A1(n4266), .A2(n4267), .ZN(n4256) );
  AOI22_X1 U3085 ( .A1(n2508), .A2(n486), .B1(n2509), .B2(n358), .ZN(n4267) );
  AOI22_X1 U3086 ( .A1(n2510), .A2(n518), .B1(n2511), .B2(n326), .ZN(n4266) );
  NAND2_X1 U3087 ( .A1(n4268), .A2(n4269), .ZN(n3202) );
  NOR4_X1 U3088 ( .A1(n4270), .A2(n4271), .A3(n4272), .A4(n4273), .ZN(n4269)
         );
  OAI21_X1 U3089 ( .B1(n1450), .B2(n2460), .A(n4274), .ZN(n4273) );
  NAND2_X1 U3090 ( .A1(n2462), .A2(n6479), .ZN(n4274) );
  OAI21_X1 U3091 ( .B1(n6103), .B2(n2463), .A(n4275), .ZN(n4272) );
  AOI22_X1 U3092 ( .A1(n2465), .A2(n6415), .B1(n2466), .B2(n6447), .ZN(n4275)
         );
  NAND2_X1 U3093 ( .A1(n4276), .A2(n4277), .ZN(n4271) );
  AOI22_X1 U3094 ( .A1(n2469), .A2(n6551), .B1(n2470), .B2(n6543), .ZN(n4277)
         );
  AOI22_X1 U3095 ( .A1(n2471), .A2(n6383), .B1(n2472), .B2(n6266), .ZN(n4276)
         );
  AOI22_X1 U3097 ( .A1(n5735), .A2(n6583), .B1(n2478), .B2(n6330), .ZN(n4281)
         );
  AOI22_X1 U3098 ( .A1(n2479), .A2(n6167), .B1(n2480), .B2(n6615), .ZN(n4280)
         );
  AOI22_X1 U3099 ( .A1(n2481), .A2(n2150), .B1(n2482), .B2(n6351), .ZN(n4279)
         );
  AOI22_X1 U3100 ( .A1(n5717), .A2(n613), .B1(n2484), .B2(n453), .ZN(n4278) );
  NOR4_X1 U3101 ( .A1(n4282), .A2(n4283), .A3(n4284), .A4(n4285), .ZN(n4268)
         );
  NAND2_X1 U3102 ( .A1(n4286), .A2(n4287), .ZN(n4285) );
  AOI22_X1 U3103 ( .A1(n2491), .A2(n389), .B1(n5709), .B2(n6199), .ZN(n4287)
         );
  AOI22_X1 U3104 ( .A1(n2493), .A2(n6298), .B1(n5457), .B2(OUT1[4]), .ZN(n4286) );
  NAND2_X1 U3105 ( .A1(n4288), .A2(n4289), .ZN(n4284) );
  AOI22_X1 U3106 ( .A1(n2496), .A2(n421), .B1(n2497), .B2(n6135), .ZN(n4289)
         );
  AOI22_X1 U3107 ( .A1(n2498), .A2(n6231), .B1(n2499), .B2(n549), .ZN(n4288)
         );
  NAND2_X1 U3108 ( .A1(n4290), .A2(n4291), .ZN(n4283) );
  AOI22_X1 U3109 ( .A1(n5691), .A2(n677), .B1(n2503), .B2(n645), .ZN(n4291) );
  AOI22_X1 U3110 ( .A1(n2504), .A2(n709), .B1(n5681), .B2(n581), .ZN(n4290) );
  NAND2_X1 U3111 ( .A1(n4292), .A2(n4293), .ZN(n4282) );
  AOI22_X1 U3112 ( .A1(n2508), .A2(n485), .B1(n2509), .B2(n357), .ZN(n4293) );
  AOI22_X1 U3113 ( .A1(n2510), .A2(n517), .B1(n2511), .B2(n325), .ZN(n4292) );
  NAND2_X1 U3114 ( .A1(n4294), .A2(n4295), .ZN(n3201) );
  NOR4_X1 U3115 ( .A1(n4296), .A2(n4297), .A3(n4298), .A4(n4299), .ZN(n4295)
         );
  OAI21_X1 U3116 ( .B1(n1451), .B2(n2460), .A(n4300), .ZN(n4299) );
  NAND2_X1 U3117 ( .A1(n2462), .A2(n6480), .ZN(n4300) );
  OAI21_X1 U3118 ( .B1(n6104), .B2(n2463), .A(n4301), .ZN(n4298) );
  AOI22_X1 U3119 ( .A1(n2465), .A2(n6416), .B1(n2466), .B2(n6448), .ZN(n4301)
         );
  NAND2_X1 U3120 ( .A1(n4302), .A2(n4303), .ZN(n4297) );
  AOI22_X1 U3121 ( .A1(n2469), .A2(n6552), .B1(n2470), .B2(n6544), .ZN(n4303)
         );
  AOI22_X1 U3122 ( .A1(n2471), .A2(n6384), .B1(n2472), .B2(n6267), .ZN(n4302)
         );
  AOI22_X1 U3124 ( .A1(n5735), .A2(n6584), .B1(n2478), .B2(n6331), .ZN(n4307)
         );
  AOI22_X1 U3125 ( .A1(n2479), .A2(n6168), .B1(n2480), .B2(n6616), .ZN(n4306)
         );
  AOI22_X1 U3126 ( .A1(n2481), .A2(n2145), .B1(n2482), .B2(n6352), .ZN(n4305)
         );
  AOI22_X1 U3127 ( .A1(n5717), .A2(n612), .B1(n2484), .B2(n452), .ZN(n4304) );
  NOR4_X1 U3128 ( .A1(n4308), .A2(n4309), .A3(n4310), .A4(n4311), .ZN(n4294)
         );
  NAND2_X1 U3129 ( .A1(n4312), .A2(n4313), .ZN(n4311) );
  AOI22_X1 U3130 ( .A1(n2491), .A2(n388), .B1(n5709), .B2(n6200), .ZN(n4313)
         );
  AOI22_X1 U3131 ( .A1(n2493), .A2(n6299), .B1(n5457), .B2(OUT1[3]), .ZN(n4312) );
  NAND2_X1 U3132 ( .A1(n4314), .A2(n4315), .ZN(n4310) );
  AOI22_X1 U3133 ( .A1(n2496), .A2(n420), .B1(n2497), .B2(n6136), .ZN(n4315)
         );
  AOI22_X1 U3134 ( .A1(n2498), .A2(n6232), .B1(n2499), .B2(n548), .ZN(n4314)
         );
  NAND2_X1 U3135 ( .A1(n4316), .A2(n4317), .ZN(n4309) );
  AOI22_X1 U3136 ( .A1(n5691), .A2(n676), .B1(n2503), .B2(n644), .ZN(n4317) );
  AOI22_X1 U3137 ( .A1(n2504), .A2(n708), .B1(n5681), .B2(n580), .ZN(n4316) );
  NAND2_X1 U3138 ( .A1(n4318), .A2(n4319), .ZN(n4308) );
  AOI22_X1 U3139 ( .A1(n2508), .A2(n484), .B1(n2509), .B2(n356), .ZN(n4319) );
  AOI22_X1 U3140 ( .A1(n2510), .A2(n516), .B1(n2511), .B2(n324), .ZN(n4318) );
  NAND2_X1 U3141 ( .A1(n4320), .A2(n4321), .ZN(n3200) );
  NOR4_X1 U3142 ( .A1(n4322), .A2(n4323), .A3(n4324), .A4(n4325), .ZN(n4321)
         );
  OAI21_X1 U3143 ( .B1(n1452), .B2(n2460), .A(n4326), .ZN(n4325) );
  NAND2_X1 U3144 ( .A1(n2462), .A2(n6481), .ZN(n4326) );
  OAI21_X1 U3145 ( .B1(n6105), .B2(n2463), .A(n4327), .ZN(n4324) );
  AOI22_X1 U3146 ( .A1(n2465), .A2(n6417), .B1(n2466), .B2(n6449), .ZN(n4327)
         );
  NAND2_X1 U3147 ( .A1(n4328), .A2(n4329), .ZN(n4323) );
  AOI22_X1 U3148 ( .A1(n2469), .A2(n6553), .B1(n2470), .B2(n6545), .ZN(n4329)
         );
  AOI22_X1 U3149 ( .A1(n2471), .A2(n6385), .B1(n2472), .B2(n6268), .ZN(n4328)
         );
  AOI22_X1 U3151 ( .A1(n5735), .A2(n6585), .B1(n2478), .B2(n6332), .ZN(n4333)
         );
  AOI22_X1 U3152 ( .A1(n2479), .A2(n6169), .B1(n2480), .B2(n6617), .ZN(n4332)
         );
  AOI22_X1 U3153 ( .A1(n2481), .A2(n2140), .B1(n2482), .B2(n6353), .ZN(n4331)
         );
  AOI22_X1 U3154 ( .A1(n5717), .A2(n611), .B1(n2484), .B2(n451), .ZN(n4330) );
  NOR4_X1 U3155 ( .A1(n4334), .A2(n4335), .A3(n4336), .A4(n4337), .ZN(n4320)
         );
  NAND2_X1 U3156 ( .A1(n4338), .A2(n4339), .ZN(n4337) );
  AOI22_X1 U3157 ( .A1(n2491), .A2(n387), .B1(n5709), .B2(n6201), .ZN(n4339)
         );
  AOI22_X1 U3158 ( .A1(n2493), .A2(n6300), .B1(n5457), .B2(OUT1[2]), .ZN(n4338) );
  NAND2_X1 U3159 ( .A1(n4340), .A2(n4341), .ZN(n4336) );
  AOI22_X1 U3160 ( .A1(n2496), .A2(n419), .B1(n2497), .B2(n6137), .ZN(n4341)
         );
  AOI22_X1 U3161 ( .A1(n2498), .A2(n6233), .B1(n2499), .B2(n547), .ZN(n4340)
         );
  NAND2_X1 U3162 ( .A1(n4342), .A2(n4343), .ZN(n4335) );
  AOI22_X1 U3163 ( .A1(n5691), .A2(n675), .B1(n2503), .B2(n643), .ZN(n4343) );
  AOI22_X1 U3164 ( .A1(n2504), .A2(n707), .B1(n5681), .B2(n579), .ZN(n4342) );
  NAND2_X1 U3165 ( .A1(n4344), .A2(n4345), .ZN(n4334) );
  AOI22_X1 U3166 ( .A1(n2508), .A2(n483), .B1(n2509), .B2(n355), .ZN(n4345) );
  AOI22_X1 U3167 ( .A1(n2510), .A2(n515), .B1(n2511), .B2(n323), .ZN(n4344) );
  NAND2_X1 U3168 ( .A1(n4346), .A2(n4347), .ZN(n3199) );
  NOR4_X1 U3169 ( .A1(n4348), .A2(n4349), .A3(n4350), .A4(n4351), .ZN(n4347)
         );
  OAI21_X1 U3170 ( .B1(n1453), .B2(n2460), .A(n4352), .ZN(n4351) );
  NAND2_X1 U3171 ( .A1(n2462), .A2(n6482), .ZN(n4352) );
  OAI21_X1 U3172 ( .B1(n6106), .B2(n2463), .A(n4353), .ZN(n4350) );
  AOI22_X1 U3173 ( .A1(n2465), .A2(n6418), .B1(n2466), .B2(n6450), .ZN(n4353)
         );
  NAND2_X1 U3174 ( .A1(n4354), .A2(n4355), .ZN(n4349) );
  AOI22_X1 U3175 ( .A1(n2469), .A2(n6554), .B1(n2470), .B2(n6546), .ZN(n4355)
         );
  AOI22_X1 U3176 ( .A1(n2471), .A2(n6386), .B1(n2472), .B2(n6269), .ZN(n4354)
         );
  AOI22_X1 U3178 ( .A1(n5735), .A2(n6586), .B1(n2478), .B2(n6333), .ZN(n4359)
         );
  AOI22_X1 U3179 ( .A1(n2479), .A2(n6170), .B1(n2480), .B2(n6618), .ZN(n4358)
         );
  AOI22_X1 U3180 ( .A1(n2481), .A2(n2135), .B1(n2482), .B2(n6354), .ZN(n4357)
         );
  AOI22_X1 U3181 ( .A1(n5717), .A2(n610), .B1(n2484), .B2(n450), .ZN(n4356) );
  NOR4_X1 U3182 ( .A1(n4360), .A2(n4361), .A3(n4362), .A4(n4363), .ZN(n4346)
         );
  NAND2_X1 U3183 ( .A1(n4364), .A2(n4365), .ZN(n4363) );
  AOI22_X1 U3184 ( .A1(n2491), .A2(n386), .B1(n5709), .B2(n6202), .ZN(n4365)
         );
  AOI22_X1 U3185 ( .A1(n5707), .A2(n6301), .B1(n5458), .B2(OUT1[1]), .ZN(n4364) );
  NAND2_X1 U3186 ( .A1(n4366), .A2(n4367), .ZN(n4362) );
  AOI22_X1 U3187 ( .A1(n2496), .A2(n418), .B1(n2497), .B2(n6138), .ZN(n4367)
         );
  AOI22_X1 U3188 ( .A1(n2498), .A2(n6234), .B1(n2499), .B2(n546), .ZN(n4366)
         );
  NAND2_X1 U3189 ( .A1(n4368), .A2(n4369), .ZN(n4361) );
  AOI22_X1 U3190 ( .A1(n5691), .A2(n674), .B1(n2503), .B2(n642), .ZN(n4369) );
  AOI22_X1 U3191 ( .A1(n2504), .A2(n706), .B1(n5681), .B2(n578), .ZN(n4368) );
  NAND2_X1 U3192 ( .A1(n4370), .A2(n4371), .ZN(n4360) );
  AOI22_X1 U3193 ( .A1(n2508), .A2(n482), .B1(n2509), .B2(n354), .ZN(n4371) );
  AOI22_X1 U3194 ( .A1(n2510), .A2(n514), .B1(n2511), .B2(n322), .ZN(n4370) );
  NAND2_X1 U3195 ( .A1(n4372), .A2(n4373), .ZN(n3198) );
  NOR4_X1 U3196 ( .A1(n4374), .A2(n4375), .A3(n4376), .A4(n4377), .ZN(n4373)
         );
  OAI21_X1 U3197 ( .B1(n1454), .B2(n2460), .A(n4378), .ZN(n4377) );
  NAND2_X1 U3198 ( .A1(n5761), .A2(n6483), .ZN(n4378) );
  NOR2_X1 U3199 ( .A1(n4379), .A2(n4380), .ZN(n2462) );
  OR2_X1 U3200 ( .A1(n4379), .A2(n4381), .ZN(n2460) );
  OAI21_X1 U3201 ( .B1(n6107), .B2(n5758), .A(n4382), .ZN(n4376) );
  AOI22_X1 U3202 ( .A1(n5755), .A2(n6419), .B1(n5752), .B2(n6451), .ZN(n4382)
         );
  NOR2_X1 U3203 ( .A1(n4381), .A2(n4383), .ZN(n2466) );
  NOR2_X1 U3204 ( .A1(n4383), .A2(n4380), .ZN(n2465) );
  NAND2_X1 U3205 ( .A1(n4384), .A2(n4385), .ZN(n2463) );
  NOR4_X1 U3206 ( .A1(n6620), .A2(n4386), .A3(n4387), .A4(n4388), .ZN(n4385)
         );
  NOR3_X1 U3207 ( .A1(n4389), .A2(n4390), .A3(n4391), .ZN(n4384) );
  NAND2_X1 U3208 ( .A1(n4392), .A2(n4393), .ZN(n4375) );
  AOI22_X1 U3209 ( .A1(n5749), .A2(n6555), .B1(n5746), .B2(n6547), .ZN(n4393)
         );
  NOR2_X1 U3210 ( .A1(n4394), .A2(n4395), .ZN(n2470) );
  NOR2_X1 U3211 ( .A1(n4395), .A2(n4396), .ZN(n2469) );
  AOI22_X1 U3212 ( .A1(n5743), .A2(n6387), .B1(n5740), .B2(n6270), .ZN(n4392)
         );
  NOR2_X1 U3213 ( .A1(n4397), .A2(n4383), .ZN(n2472) );
  NOR2_X1 U3214 ( .A1(n4395), .A2(n4381), .ZN(n2471) );
  AOI22_X1 U3216 ( .A1(n5735), .A2(n6587), .B1(n5734), .B2(n6334), .ZN(n4401)
         );
  NOR2_X1 U3217 ( .A1(n4402), .A2(n4379), .ZN(n2478) );
  NOR2_X1 U3218 ( .A1(n4403), .A2(n4394), .ZN(n2477) );
  AOI22_X1 U3219 ( .A1(n5731), .A2(n6171), .B1(n5728), .B2(n6619), .ZN(n4400)
         );
  NOR2_X1 U3220 ( .A1(n4403), .A2(n4396), .ZN(n2480) );
  NOR2_X1 U3221 ( .A1(n4403), .A2(n4404), .ZN(n2479) );
  AOI22_X1 U3222 ( .A1(n5725), .A2(n2130), .B1(n5722), .B2(n6355), .ZN(n4399)
         );
  NOR2_X1 U3223 ( .A1(n4397), .A2(n4379), .ZN(n2482) );
  NOR2_X1 U3224 ( .A1(n4402), .A2(n4383), .ZN(n2481) );
  AOI22_X1 U3225 ( .A1(n5717), .A2(n609), .B1(n5716), .B2(n449), .ZN(n4398) );
  NOR2_X1 U3226 ( .A1(n4405), .A2(n4379), .ZN(n2484) );
  NOR2_X1 U3227 ( .A1(n4405), .A2(n4395), .ZN(n2483) );
  NOR4_X1 U3228 ( .A1(n4406), .A2(n4407), .A3(n4408), .A4(n4409), .ZN(n4372)
         );
  NAND2_X1 U3229 ( .A1(n4410), .A2(n4411), .ZN(n4409) );
  AOI22_X1 U3230 ( .A1(n5713), .A2(n385), .B1(n5709), .B2(n6203), .ZN(n4411)
         );
  NOR2_X1 U3231 ( .A1(n4405), .A2(n4403), .ZN(n2492) );
  NOR2_X1 U3232 ( .A1(n4402), .A2(n4403), .ZN(n2491) );
  AOI22_X1 U3233 ( .A1(n5707), .A2(n6302), .B1(n5458), .B2(OUT1[0]), .ZN(n4410) );
  NOR2_X1 U3234 ( .A1(n4403), .A2(n4397), .ZN(n2493) );
  NAND2_X1 U3235 ( .A1(n4412), .A2(n4413), .ZN(n4408) );
  AOI22_X1 U3236 ( .A1(n5704), .A2(n417), .B1(n5701), .B2(n6139), .ZN(n4413)
         );
  NOR2_X1 U3237 ( .A1(n4383), .A2(n4404), .ZN(n2497) );
  NOR2_X1 U3238 ( .A1(n4397), .A2(n4395), .ZN(n2496) );
  NAND2_X1 U3239 ( .A1(n4414), .A2(ADD_RD1[3]), .ZN(n4397) );
  NOR2_X1 U3240 ( .A1(ADD_RD1[4]), .A2(n6071), .ZN(n4414) );
  AOI22_X1 U3241 ( .A1(n5698), .A2(n6235), .B1(n5695), .B2(n545), .ZN(n4412)
         );
  NOR2_X1 U3242 ( .A1(n4402), .A2(n4395), .ZN(n2499) );
  NAND2_X1 U3243 ( .A1(n4415), .A2(ADD_RD1[3]), .ZN(n4402) );
  NOR2_X1 U3244 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[0]), .ZN(n4415) );
  NOR2_X1 U3245 ( .A1(n4379), .A2(n4404), .ZN(n2498) );
  NAND2_X1 U3246 ( .A1(n4416), .A2(n4417), .ZN(n4407) );
  AOI22_X1 U3247 ( .A1(n2502), .A2(n673), .B1(n5689), .B2(n641), .ZN(n4417) );
  NOR2_X1 U3248 ( .A1(n4396), .A2(n4383), .ZN(n2503) );
  NOR2_X1 U3249 ( .A1(n4395), .A2(n4380), .ZN(n2502) );
  NAND2_X1 U3250 ( .A1(n4418), .A2(n4419), .ZN(n4395) );
  NOR2_X1 U3251 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n4418) );
  AOI22_X1 U3252 ( .A1(n5686), .A2(n705), .B1(n5681), .B2(n577), .ZN(n4416) );
  NOR2_X1 U3253 ( .A1(n4405), .A2(n4383), .ZN(n2505) );
  OR2_X1 U3254 ( .A1(n4420), .A2(n6071), .ZN(n4405) );
  OR2_X1 U3255 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n4420) );
  NOR2_X1 U3256 ( .A1(n4403), .A2(n4380), .ZN(n2504) );
  OR2_X1 U3257 ( .A1(n4421), .A2(n6068), .ZN(n4380) );
  OR2_X1 U3258 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .ZN(n4421) );
  NAND2_X1 U3259 ( .A1(n4422), .A2(n4423), .ZN(n4406) );
  AOI22_X1 U3260 ( .A1(n5680), .A2(n481), .B1(n5677), .B2(n353), .ZN(n4423) );
  NOR2_X1 U3261 ( .A1(n4394), .A2(n4379), .ZN(n2509) );
  NOR2_X1 U3262 ( .A1(n4394), .A2(n4383), .ZN(n2508) );
  NAND2_X1 U3263 ( .A1(n4424), .A2(n4419), .ZN(n4383) );
  NOR2_X1 U3264 ( .A1(ADD_RD1[2]), .A2(n6070), .ZN(n4424) );
  NAND2_X1 U3265 ( .A1(n4425), .A2(ADD_RD1[3]), .ZN(n4394) );
  NOR2_X1 U3266 ( .A1(ADD_RD1[0]), .A2(n6068), .ZN(n4425) );
  AOI22_X1 U3267 ( .A1(n5674), .A2(n513), .B1(n5671), .B2(n321), .ZN(n4422) );
  NOR2_X1 U3268 ( .A1(n4396), .A2(n4379), .ZN(n2511) );
  NAND2_X1 U3269 ( .A1(n4426), .A2(n4419), .ZN(n4379) );
  NOR2_X1 U3270 ( .A1(n6069), .A2(n6070), .ZN(n4426) );
  NAND2_X1 U3271 ( .A1(n4427), .A2(ADD_RD1[3]), .ZN(n4396) );
  NOR2_X1 U3272 ( .A1(n6068), .A2(n6071), .ZN(n4427) );
  NOR2_X1 U3273 ( .A1(n4403), .A2(n4381), .ZN(n2510) );
  OR2_X1 U3274 ( .A1(n4428), .A2(n6071), .ZN(n4381) );
  OR2_X1 U3275 ( .A1(ADD_RD1[3]), .A2(n6068), .ZN(n4428) );
  NAND2_X1 U3276 ( .A1(n4429), .A2(n4419), .ZN(n4403) );
  NOR2_X1 U3277 ( .A1(n4389), .A2(n4430), .ZN(n4419) );
  XOR2_X1 U3280 ( .A(ADD_WR[3]), .B(ADD_RD1[3]), .Z(n4386) );
  XOR2_X1 U3281 ( .A(ADD_RD1[1]), .B(ADD_WR[1]), .Z(n4387) );
  XOR2_X1 U3283 ( .A(ADD_WR[4]), .B(ADD_RD1[4]), .Z(n4390) );
  XOR2_X1 U3284 ( .A(ADD_RD1[0]), .B(ADD_WR[0]), .Z(n4388) );
  XOR2_X1 U3285 ( .A(ADD_RD1[2]), .B(ADD_WR[2]), .Z(n4391) );
  NAND2_X1 U3286 ( .A1(n4433), .A2(RD1), .ZN(n4389) );
  NOR2_X1 U3287 ( .A1(n4434), .A2(n5939), .ZN(n4433) );
  NOR3_X1 U3288 ( .A1(n4404), .A2(ADD_RD1[2]), .A3(ADD_RD1[1]), .ZN(n4434) );
  NAND2_X1 U3289 ( .A1(n4435), .A2(n6071), .ZN(n4404) );
  NOR2_X1 U3290 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n4435) );
  NOR2_X1 U3291 ( .A1(ADD_RD1[1]), .A2(n6069), .ZN(n4429) );
  NAND2_X1 U3292 ( .A1(n4436), .A2(n4437), .ZN(n3197) );
  NOR4_X1 U3293 ( .A1(n4438), .A2(n4439), .A3(n4440), .A4(n4441), .ZN(n4437)
         );
  OAI21_X1 U3294 ( .B1(n1423), .B2(n5668), .A(n4443), .ZN(n4441) );
  NAND2_X1 U3295 ( .A1(n4444), .A2(n6452), .ZN(n4443) );
  OAI21_X1 U3296 ( .B1(n6076), .B2(n5662), .A(n4446), .ZN(n4440) );
  AOI22_X1 U3297 ( .A1(n5659), .A2(n6388), .B1(n5656), .B2(n6420), .ZN(n4446)
         );
  NAND2_X1 U3298 ( .A1(n4449), .A2(n4450), .ZN(n4439) );
  AOI22_X1 U3299 ( .A1(n5653), .A2(n2830), .B1(n5650), .B2(n6516), .ZN(n4450)
         );
  AOI22_X1 U3300 ( .A1(n5645), .A2(n6356), .B1(n5644), .B2(n6556), .ZN(n4449)
         );
  AOI22_X1 U3302 ( .A1(n5641), .A2(n2382), .B1(n5638), .B2(n6303), .ZN(n4458)
         );
  AOI22_X1 U3303 ( .A1(n5634), .A2(n6140), .B1(n5632), .B2(n6588), .ZN(n4457)
         );
  AOI22_X1 U3304 ( .A1(n5629), .A2(n6236), .B1(n5626), .B2(n6239), .ZN(n4456)
         );
  AOI22_X1 U3305 ( .A1(n5623), .A2(n640), .B1(n5620), .B2(n480), .ZN(n4455) );
  NOR4_X1 U3306 ( .A1(n4467), .A2(n4468), .A3(n4469), .A4(n4470), .ZN(n4436)
         );
  NAND2_X1 U3307 ( .A1(n4471), .A2(n4472), .ZN(n4470) );
  AOI22_X1 U3308 ( .A1(n5617), .A2(n416), .B1(n5614), .B2(n6172), .ZN(n4472)
         );
  AOI22_X1 U3309 ( .A1(n5611), .A2(n6271), .B1(n5458), .B2(OUT2[31]), .ZN(
        n4471) );
  NAND2_X1 U3310 ( .A1(n4476), .A2(n4477), .ZN(n4469) );
  AOI22_X1 U3311 ( .A1(n5608), .A2(n448), .B1(n5605), .B2(n6108), .ZN(n4477)
         );
  AOI22_X1 U3312 ( .A1(n5602), .A2(n6204), .B1(n4481), .B2(n576), .ZN(n4476)
         );
  NAND2_X1 U3313 ( .A1(n4482), .A2(n4483), .ZN(n4468) );
  AOI22_X1 U3314 ( .A1(n5596), .A2(n704), .B1(n5591), .B2(n672), .ZN(n4483) );
  AOI22_X1 U3315 ( .A1(n5590), .A2(n736), .B1(n5587), .B2(n608), .ZN(n4482) );
  NAND2_X1 U3316 ( .A1(n4488), .A2(n4489), .ZN(n4467) );
  AOI22_X1 U3317 ( .A1(n5584), .A2(n512), .B1(n5581), .B2(n384), .ZN(n4489) );
  AOI22_X1 U3318 ( .A1(n5578), .A2(n544), .B1(n5573), .B2(n352), .ZN(n4488) );
  NAND2_X1 U3319 ( .A1(n4494), .A2(n4495), .ZN(n3196) );
  NOR4_X1 U3320 ( .A1(n4496), .A2(n4497), .A3(n4498), .A4(n4499), .ZN(n4495)
         );
  OAI21_X1 U3321 ( .B1(n1424), .B2(n5668), .A(n4500), .ZN(n4499) );
  NAND2_X1 U3322 ( .A1(n4444), .A2(n6453), .ZN(n4500) );
  OAI21_X1 U3323 ( .B1(n6077), .B2(n5662), .A(n4501), .ZN(n4498) );
  AOI22_X1 U3324 ( .A1(n5659), .A2(n6389), .B1(n5656), .B2(n6421), .ZN(n4501)
         );
  NAND2_X1 U3325 ( .A1(n4502), .A2(n4503), .ZN(n4497) );
  AOI22_X1 U3326 ( .A1(n5653), .A2(n2829), .B1(n5650), .B2(n6517), .ZN(n4503)
         );
  AOI22_X1 U3327 ( .A1(n5645), .A2(n6357), .B1(n5644), .B2(n6557), .ZN(n4502)
         );
  AOI22_X1 U3329 ( .A1(n5641), .A2(n2379), .B1(n5638), .B2(n6304), .ZN(n4507)
         );
  AOI22_X1 U3330 ( .A1(n4461), .A2(n6141), .B1(n5632), .B2(n6589), .ZN(n4506)
         );
  AOI22_X1 U3331 ( .A1(n5629), .A2(n6237), .B1(n5626), .B2(n6240), .ZN(n4505)
         );
  AOI22_X1 U3332 ( .A1(n5623), .A2(n639), .B1(n5620), .B2(n479), .ZN(n4504) );
  NOR4_X1 U3333 ( .A1(n4508), .A2(n4509), .A3(n4510), .A4(n4511), .ZN(n4494)
         );
  NAND2_X1 U3334 ( .A1(n4512), .A2(n4513), .ZN(n4511) );
  AOI22_X1 U3335 ( .A1(n5617), .A2(n415), .B1(n5614), .B2(n6173), .ZN(n4513)
         );
  AOI22_X1 U3336 ( .A1(n5611), .A2(n6272), .B1(n5457), .B2(OUT2[30]), .ZN(
        n4512) );
  NAND2_X1 U3337 ( .A1(n4514), .A2(n4515), .ZN(n4510) );
  AOI22_X1 U3338 ( .A1(n5608), .A2(n447), .B1(n5605), .B2(n6109), .ZN(n4515)
         );
  AOI22_X1 U3339 ( .A1(n5602), .A2(n6205), .B1(n4481), .B2(n575), .ZN(n4514)
         );
  NAND2_X1 U3340 ( .A1(n4516), .A2(n4517), .ZN(n4509) );
  AOI22_X1 U3341 ( .A1(n5596), .A2(n703), .B1(n5591), .B2(n671), .ZN(n4517) );
  AOI22_X1 U3342 ( .A1(n5590), .A2(n735), .B1(n5587), .B2(n607), .ZN(n4516) );
  NAND2_X1 U3343 ( .A1(n4518), .A2(n4519), .ZN(n4508) );
  AOI22_X1 U3344 ( .A1(n5584), .A2(n511), .B1(n5581), .B2(n383), .ZN(n4519) );
  AOI22_X1 U3345 ( .A1(n5578), .A2(n543), .B1(n5573), .B2(n351), .ZN(n4518) );
  NAND2_X1 U3346 ( .A1(n4520), .A2(n4521), .ZN(n3195) );
  NOR4_X1 U3347 ( .A1(n4522), .A2(n4523), .A3(n4524), .A4(n4525), .ZN(n4521)
         );
  OAI21_X1 U3348 ( .B1(n1425), .B2(n5668), .A(n4526), .ZN(n4525) );
  NAND2_X1 U3349 ( .A1(n4444), .A2(n6454), .ZN(n4526) );
  OAI21_X1 U3350 ( .B1(n6078), .B2(n5662), .A(n4527), .ZN(n4524) );
  AOI22_X1 U3351 ( .A1(n5659), .A2(n6390), .B1(n5656), .B2(n6422), .ZN(n4527)
         );
  NAND2_X1 U3352 ( .A1(n4528), .A2(n4529), .ZN(n4523) );
  AOI22_X1 U3353 ( .A1(n5653), .A2(n2828), .B1(n5650), .B2(n6518), .ZN(n4529)
         );
  AOI22_X1 U3354 ( .A1(n5645), .A2(n6358), .B1(n5644), .B2(n6558), .ZN(n4528)
         );
  AOI22_X1 U3356 ( .A1(n5641), .A2(n2376), .B1(n5638), .B2(n6305), .ZN(n4533)
         );
  AOI22_X1 U3357 ( .A1(n4461), .A2(n6142), .B1(n5632), .B2(n6590), .ZN(n4532)
         );
  AOI22_X1 U3358 ( .A1(n5629), .A2(n6238), .B1(n5626), .B2(n6241), .ZN(n4531)
         );
  AOI22_X1 U3359 ( .A1(n5623), .A2(n638), .B1(n5620), .B2(n478), .ZN(n4530) );
  NOR4_X1 U3360 ( .A1(n4534), .A2(n4535), .A3(n4536), .A4(n4537), .ZN(n4520)
         );
  NAND2_X1 U3361 ( .A1(n4538), .A2(n4539), .ZN(n4537) );
  AOI22_X1 U3362 ( .A1(n5617), .A2(n414), .B1(n5614), .B2(n6174), .ZN(n4539)
         );
  AOI22_X1 U3363 ( .A1(n5611), .A2(n6273), .B1(n5457), .B2(OUT2[29]), .ZN(
        n4538) );
  NAND2_X1 U3364 ( .A1(n4540), .A2(n4541), .ZN(n4536) );
  AOI22_X1 U3365 ( .A1(n5608), .A2(n446), .B1(n5605), .B2(n6110), .ZN(n4541)
         );
  AOI22_X1 U3366 ( .A1(n5602), .A2(n6206), .B1(n4481), .B2(n574), .ZN(n4540)
         );
  NAND2_X1 U3367 ( .A1(n4542), .A2(n4543), .ZN(n4535) );
  AOI22_X1 U3368 ( .A1(n5596), .A2(n702), .B1(n5591), .B2(n670), .ZN(n4543) );
  AOI22_X1 U3369 ( .A1(n5590), .A2(n734), .B1(n5587), .B2(n606), .ZN(n4542) );
  NAND2_X1 U3370 ( .A1(n4544), .A2(n4545), .ZN(n4534) );
  AOI22_X1 U3371 ( .A1(n5584), .A2(n510), .B1(n5581), .B2(n382), .ZN(n4545) );
  AOI22_X1 U3372 ( .A1(n5578), .A2(n542), .B1(n5573), .B2(n350), .ZN(n4544) );
  NAND2_X1 U3373 ( .A1(n4546), .A2(n4547), .ZN(n3194) );
  NOR4_X1 U3374 ( .A1(n4548), .A2(n4549), .A3(n4550), .A4(n4551), .ZN(n4547)
         );
  OAI21_X1 U3375 ( .B1(n1426), .B2(n5668), .A(n4552), .ZN(n4551) );
  NAND2_X1 U3376 ( .A1(n4444), .A2(n6455), .ZN(n4552) );
  OAI21_X1 U3377 ( .B1(n6079), .B2(n5662), .A(n4553), .ZN(n4550) );
  AOI22_X1 U3378 ( .A1(n5659), .A2(n6391), .B1(n5656), .B2(n6423), .ZN(n4553)
         );
  NAND2_X1 U3379 ( .A1(n4554), .A2(n4555), .ZN(n4549) );
  AOI22_X1 U3380 ( .A1(n5653), .A2(n2827), .B1(n5650), .B2(n6519), .ZN(n4555)
         );
  AOI22_X1 U3381 ( .A1(n5645), .A2(n6359), .B1(n5644), .B2(n6559), .ZN(n4554)
         );
  AOI22_X1 U3383 ( .A1(n5641), .A2(n2373), .B1(n5638), .B2(n6306), .ZN(n4559)
         );
  AOI22_X1 U3384 ( .A1(n4461), .A2(n6143), .B1(n5632), .B2(n6591), .ZN(n4558)
         );
  AOI22_X1 U3385 ( .A1(n5629), .A2(n2270), .B1(n5626), .B2(n6242), .ZN(n4557)
         );
  AOI22_X1 U3386 ( .A1(n5623), .A2(n637), .B1(n5620), .B2(n477), .ZN(n4556) );
  NOR4_X1 U3387 ( .A1(n4560), .A2(n4561), .A3(n4562), .A4(n4563), .ZN(n4546)
         );
  NAND2_X1 U3388 ( .A1(n4564), .A2(n4565), .ZN(n4563) );
  AOI22_X1 U3389 ( .A1(n5617), .A2(n413), .B1(n5614), .B2(n6175), .ZN(n4565)
         );
  AOI22_X1 U3390 ( .A1(n5611), .A2(n6274), .B1(n5457), .B2(OUT2[28]), .ZN(
        n4564) );
  NAND2_X1 U3391 ( .A1(n4566), .A2(n4567), .ZN(n4562) );
  AOI22_X1 U3392 ( .A1(n5608), .A2(n445), .B1(n5605), .B2(n6111), .ZN(n4567)
         );
  AOI22_X1 U3393 ( .A1(n5602), .A2(n6207), .B1(n4481), .B2(n573), .ZN(n4566)
         );
  NAND2_X1 U3394 ( .A1(n4568), .A2(n4569), .ZN(n4561) );
  AOI22_X1 U3395 ( .A1(n5596), .A2(n701), .B1(n5591), .B2(n669), .ZN(n4569) );
  AOI22_X1 U3396 ( .A1(n5590), .A2(n733), .B1(n5587), .B2(n605), .ZN(n4568) );
  NAND2_X1 U3397 ( .A1(n4570), .A2(n4571), .ZN(n4560) );
  AOI22_X1 U3398 ( .A1(n5584), .A2(n509), .B1(n5581), .B2(n381), .ZN(n4571) );
  AOI22_X1 U3399 ( .A1(n5578), .A2(n541), .B1(n5573), .B2(n349), .ZN(n4570) );
  NAND2_X1 U3400 ( .A1(n4572), .A2(n4573), .ZN(n3193) );
  NOR4_X1 U3401 ( .A1(n4574), .A2(n4575), .A3(n4576), .A4(n4577), .ZN(n4573)
         );
  OAI21_X1 U3402 ( .B1(n1427), .B2(n5668), .A(n4578), .ZN(n4577) );
  NAND2_X1 U3403 ( .A1(n4444), .A2(n6456), .ZN(n4578) );
  OAI21_X1 U3404 ( .B1(n6080), .B2(n5662), .A(n4579), .ZN(n4576) );
  AOI22_X1 U3405 ( .A1(n5659), .A2(n6392), .B1(n5656), .B2(n6424), .ZN(n4579)
         );
  NAND2_X1 U3406 ( .A1(n4580), .A2(n4581), .ZN(n4575) );
  AOI22_X1 U3407 ( .A1(n5653), .A2(n2826), .B1(n5650), .B2(n6520), .ZN(n4581)
         );
  AOI22_X1 U3408 ( .A1(n5645), .A2(n6360), .B1(n5644), .B2(n6560), .ZN(n4580)
         );
  AOI22_X1 U3410 ( .A1(n5641), .A2(n2370), .B1(n5638), .B2(n6307), .ZN(n4585)
         );
  AOI22_X1 U3411 ( .A1(n4461), .A2(n6144), .B1(n5632), .B2(n6592), .ZN(n4584)
         );
  AOI22_X1 U3412 ( .A1(n5629), .A2(n2265), .B1(n5626), .B2(n6243), .ZN(n4583)
         );
  AOI22_X1 U3413 ( .A1(n5623), .A2(n636), .B1(n5620), .B2(n476), .ZN(n4582) );
  NOR4_X1 U3414 ( .A1(n4586), .A2(n4587), .A3(n4588), .A4(n4589), .ZN(n4572)
         );
  NAND2_X1 U3415 ( .A1(n4590), .A2(n4591), .ZN(n4589) );
  AOI22_X1 U3416 ( .A1(n5617), .A2(n412), .B1(n5614), .B2(n6176), .ZN(n4591)
         );
  AOI22_X1 U3417 ( .A1(n5611), .A2(n6275), .B1(n5457), .B2(OUT2[27]), .ZN(
        n4590) );
  NAND2_X1 U3418 ( .A1(n4592), .A2(n4593), .ZN(n4588) );
  AOI22_X1 U3419 ( .A1(n5608), .A2(n444), .B1(n5605), .B2(n6112), .ZN(n4593)
         );
  AOI22_X1 U3420 ( .A1(n5602), .A2(n6208), .B1(n4481), .B2(n572), .ZN(n4592)
         );
  NAND2_X1 U3421 ( .A1(n4594), .A2(n4595), .ZN(n4587) );
  AOI22_X1 U3422 ( .A1(n5596), .A2(n700), .B1(n5591), .B2(n668), .ZN(n4595) );
  AOI22_X1 U3423 ( .A1(n5590), .A2(n732), .B1(n5587), .B2(n604), .ZN(n4594) );
  NAND2_X1 U3424 ( .A1(n4596), .A2(n4597), .ZN(n4586) );
  AOI22_X1 U3425 ( .A1(n5584), .A2(n508), .B1(n5581), .B2(n380), .ZN(n4597) );
  AOI22_X1 U3426 ( .A1(n5578), .A2(n540), .B1(n5573), .B2(n348), .ZN(n4596) );
  NAND2_X1 U3427 ( .A1(n4598), .A2(n4599), .ZN(n3192) );
  NOR4_X1 U3428 ( .A1(n4600), .A2(n4601), .A3(n4602), .A4(n4603), .ZN(n4599)
         );
  OAI21_X1 U3429 ( .B1(n1428), .B2(n5668), .A(n4604), .ZN(n4603) );
  NAND2_X1 U3430 ( .A1(n4444), .A2(n6457), .ZN(n4604) );
  OAI21_X1 U3431 ( .B1(n6081), .B2(n5662), .A(n4605), .ZN(n4602) );
  AOI22_X1 U3432 ( .A1(n5659), .A2(n6393), .B1(n5656), .B2(n6425), .ZN(n4605)
         );
  NAND2_X1 U3433 ( .A1(n4606), .A2(n4607), .ZN(n4601) );
  AOI22_X1 U3434 ( .A1(n5653), .A2(n2825), .B1(n5650), .B2(n6521), .ZN(n4607)
         );
  AOI22_X1 U3435 ( .A1(n5645), .A2(n6361), .B1(n5644), .B2(n6561), .ZN(n4606)
         );
  AOI22_X1 U3437 ( .A1(n5641), .A2(n2367), .B1(n5638), .B2(n6308), .ZN(n4611)
         );
  AOI22_X1 U3438 ( .A1(n4461), .A2(n6145), .B1(n5632), .B2(n6593), .ZN(n4610)
         );
  AOI22_X1 U3439 ( .A1(n5629), .A2(n2260), .B1(n5626), .B2(n6244), .ZN(n4609)
         );
  AOI22_X1 U3440 ( .A1(n5623), .A2(n635), .B1(n5620), .B2(n475), .ZN(n4608) );
  NOR4_X1 U3441 ( .A1(n4612), .A2(n4613), .A3(n4614), .A4(n4615), .ZN(n4598)
         );
  NAND2_X1 U3442 ( .A1(n4616), .A2(n4617), .ZN(n4615) );
  AOI22_X1 U3443 ( .A1(n5617), .A2(n411), .B1(n5614), .B2(n6177), .ZN(n4617)
         );
  AOI22_X1 U3444 ( .A1(n5611), .A2(n6276), .B1(n5457), .B2(OUT2[26]), .ZN(
        n4616) );
  NAND2_X1 U3445 ( .A1(n4618), .A2(n4619), .ZN(n4614) );
  AOI22_X1 U3446 ( .A1(n5608), .A2(n443), .B1(n5605), .B2(n6113), .ZN(n4619)
         );
  AOI22_X1 U3447 ( .A1(n5602), .A2(n6209), .B1(n4481), .B2(n571), .ZN(n4618)
         );
  NAND2_X1 U3448 ( .A1(n4620), .A2(n4621), .ZN(n4613) );
  AOI22_X1 U3449 ( .A1(n5596), .A2(n699), .B1(n5591), .B2(n667), .ZN(n4621) );
  AOI22_X1 U3450 ( .A1(n5590), .A2(n731), .B1(n5587), .B2(n603), .ZN(n4620) );
  NAND2_X1 U3451 ( .A1(n4622), .A2(n4623), .ZN(n4612) );
  AOI22_X1 U3452 ( .A1(n5584), .A2(n507), .B1(n5581), .B2(n379), .ZN(n4623) );
  AOI22_X1 U3453 ( .A1(n5578), .A2(n539), .B1(n5573), .B2(n347), .ZN(n4622) );
  NAND2_X1 U3454 ( .A1(n4624), .A2(n4625), .ZN(n3191) );
  NOR4_X1 U3455 ( .A1(n4626), .A2(n4627), .A3(n4628), .A4(n4629), .ZN(n4625)
         );
  OAI21_X1 U3456 ( .B1(n1429), .B2(n5668), .A(n4630), .ZN(n4629) );
  NAND2_X1 U3457 ( .A1(n4444), .A2(n6458), .ZN(n4630) );
  OAI21_X1 U3458 ( .B1(n5477), .B2(n5662), .A(n4631), .ZN(n4628) );
  AOI22_X1 U3459 ( .A1(n5659), .A2(n6394), .B1(n5656), .B2(n6426), .ZN(n4631)
         );
  NAND2_X1 U3460 ( .A1(n4632), .A2(n4633), .ZN(n4627) );
  AOI22_X1 U3461 ( .A1(n5653), .A2(n2824), .B1(n5650), .B2(n6522), .ZN(n4633)
         );
  AOI22_X1 U3462 ( .A1(n5645), .A2(n6362), .B1(n5644), .B2(n6562), .ZN(n4632)
         );
  AOI22_X1 U3464 ( .A1(n5641), .A2(n2364), .B1(n5638), .B2(n6309), .ZN(n4637)
         );
  AOI22_X1 U3465 ( .A1(n4461), .A2(n6146), .B1(n5632), .B2(n6594), .ZN(n4636)
         );
  AOI22_X1 U3466 ( .A1(n5629), .A2(n2255), .B1(n5626), .B2(n6245), .ZN(n4635)
         );
  AOI22_X1 U3467 ( .A1(n5623), .A2(n634), .B1(n5620), .B2(n474), .ZN(n4634) );
  NOR4_X1 U3468 ( .A1(n4638), .A2(n4639), .A3(n4640), .A4(n4641), .ZN(n4624)
         );
  NAND2_X1 U3469 ( .A1(n4642), .A2(n4643), .ZN(n4641) );
  AOI22_X1 U3470 ( .A1(n5617), .A2(n410), .B1(n5614), .B2(n6178), .ZN(n4643)
         );
  AOI22_X1 U3471 ( .A1(n5611), .A2(n6277), .B1(n5457), .B2(OUT2[25]), .ZN(
        n4642) );
  NAND2_X1 U3472 ( .A1(n4644), .A2(n4645), .ZN(n4640) );
  AOI22_X1 U3473 ( .A1(n5608), .A2(n442), .B1(n5605), .B2(n6114), .ZN(n4645)
         );
  AOI22_X1 U3474 ( .A1(n5602), .A2(n6210), .B1(n4481), .B2(n570), .ZN(n4644)
         );
  NAND2_X1 U3475 ( .A1(n4646), .A2(n4647), .ZN(n4639) );
  AOI22_X1 U3476 ( .A1(n5596), .A2(n698), .B1(n5591), .B2(n666), .ZN(n4647) );
  AOI22_X1 U3477 ( .A1(n5590), .A2(n730), .B1(n5587), .B2(n602), .ZN(n4646) );
  NAND2_X1 U3478 ( .A1(n4648), .A2(n4649), .ZN(n4638) );
  AOI22_X1 U3479 ( .A1(n5584), .A2(n506), .B1(n5581), .B2(n378), .ZN(n4649) );
  AOI22_X1 U3480 ( .A1(n5578), .A2(n538), .B1(n5573), .B2(n346), .ZN(n4648) );
  NAND2_X1 U3481 ( .A1(n4650), .A2(n4651), .ZN(n3190) );
  NOR4_X1 U3482 ( .A1(n4652), .A2(n4653), .A3(n4654), .A4(n4655), .ZN(n4651)
         );
  OAI21_X1 U3483 ( .B1(n1430), .B2(n5668), .A(n4656), .ZN(n4655) );
  NAND2_X1 U3484 ( .A1(n4444), .A2(n6459), .ZN(n4656) );
  OAI21_X1 U3485 ( .B1(n6083), .B2(n5662), .A(n4657), .ZN(n4654) );
  AOI22_X1 U3486 ( .A1(n5659), .A2(n6395), .B1(n5656), .B2(n6427), .ZN(n4657)
         );
  NAND2_X1 U3487 ( .A1(n4658), .A2(n4659), .ZN(n4653) );
  AOI22_X1 U3488 ( .A1(n5653), .A2(n2823), .B1(n5650), .B2(n6523), .ZN(n4659)
         );
  AOI22_X1 U3489 ( .A1(n5645), .A2(n6363), .B1(n5644), .B2(n6563), .ZN(n4658)
         );
  AOI22_X1 U3491 ( .A1(n5641), .A2(n2361), .B1(n5638), .B2(n6310), .ZN(n4663)
         );
  AOI22_X1 U3492 ( .A1(n4461), .A2(n6147), .B1(n5632), .B2(n6595), .ZN(n4662)
         );
  AOI22_X1 U3493 ( .A1(n5629), .A2(n2250), .B1(n5626), .B2(n6246), .ZN(n4661)
         );
  AOI22_X1 U3494 ( .A1(n5623), .A2(n633), .B1(n5620), .B2(n473), .ZN(n4660) );
  NOR4_X1 U3495 ( .A1(n4664), .A2(n4665), .A3(n4666), .A4(n4667), .ZN(n4650)
         );
  NAND2_X1 U3496 ( .A1(n4668), .A2(n4669), .ZN(n4667) );
  AOI22_X1 U3497 ( .A1(n5617), .A2(n409), .B1(n5614), .B2(n6179), .ZN(n4669)
         );
  AOI22_X1 U3498 ( .A1(n5611), .A2(n6278), .B1(n5457), .B2(OUT2[24]), .ZN(
        n4668) );
  NAND2_X1 U3499 ( .A1(n4670), .A2(n4671), .ZN(n4666) );
  AOI22_X1 U3500 ( .A1(n5608), .A2(n441), .B1(n5605), .B2(n6115), .ZN(n4671)
         );
  AOI22_X1 U3501 ( .A1(n5602), .A2(n6211), .B1(n4481), .B2(n569), .ZN(n4670)
         );
  NAND2_X1 U3502 ( .A1(n4672), .A2(n4673), .ZN(n4665) );
  AOI22_X1 U3503 ( .A1(n5596), .A2(n697), .B1(n5591), .B2(n665), .ZN(n4673) );
  AOI22_X1 U3504 ( .A1(n5590), .A2(n729), .B1(n5587), .B2(n601), .ZN(n4672) );
  NAND2_X1 U3505 ( .A1(n4674), .A2(n4675), .ZN(n4664) );
  AOI22_X1 U3506 ( .A1(n5584), .A2(n505), .B1(n5581), .B2(n377), .ZN(n4675) );
  AOI22_X1 U3507 ( .A1(n5578), .A2(n537), .B1(n5573), .B2(n345), .ZN(n4674) );
  NAND2_X1 U3508 ( .A1(n4676), .A2(n4677), .ZN(n3189) );
  NOR4_X1 U3509 ( .A1(n4678), .A2(n4679), .A3(n4680), .A4(n4681), .ZN(n4677)
         );
  OAI21_X1 U3510 ( .B1(n1431), .B2(n5668), .A(n4682), .ZN(n4681) );
  NAND2_X1 U3511 ( .A1(n4444), .A2(n6460), .ZN(n4682) );
  OAI21_X1 U3512 ( .B1(n6084), .B2(n5662), .A(n4683), .ZN(n4680) );
  AOI22_X1 U3513 ( .A1(n5659), .A2(n6396), .B1(n5656), .B2(n6428), .ZN(n4683)
         );
  NAND2_X1 U3514 ( .A1(n4684), .A2(n4685), .ZN(n4679) );
  AOI22_X1 U3515 ( .A1(n5653), .A2(n2822), .B1(n5650), .B2(n6524), .ZN(n4685)
         );
  AOI22_X1 U3516 ( .A1(n4453), .A2(n6364), .B1(n5644), .B2(n6564), .ZN(n4684)
         );
  AOI22_X1 U3518 ( .A1(n5641), .A2(n2358), .B1(n5638), .B2(n6311), .ZN(n4689)
         );
  AOI22_X1 U3519 ( .A1(n4461), .A2(n6148), .B1(n5632), .B2(n6596), .ZN(n4688)
         );
  AOI22_X1 U3520 ( .A1(n5629), .A2(n2245), .B1(n5626), .B2(n6247), .ZN(n4687)
         );
  AOI22_X1 U3521 ( .A1(n5623), .A2(n632), .B1(n5620), .B2(n472), .ZN(n4686) );
  NOR4_X1 U3522 ( .A1(n4690), .A2(n4691), .A3(n4692), .A4(n4693), .ZN(n4676)
         );
  NAND2_X1 U3523 ( .A1(n4694), .A2(n4695), .ZN(n4693) );
  AOI22_X1 U3524 ( .A1(n5617), .A2(n408), .B1(n5614), .B2(n6180), .ZN(n4695)
         );
  AOI22_X1 U3525 ( .A1(n5611), .A2(n6279), .B1(n5457), .B2(OUT2[23]), .ZN(
        n4694) );
  NAND2_X1 U3526 ( .A1(n4696), .A2(n4697), .ZN(n4692) );
  AOI22_X1 U3527 ( .A1(n5608), .A2(n440), .B1(n5605), .B2(n6116), .ZN(n4697)
         );
  AOI22_X1 U3528 ( .A1(n5602), .A2(n6212), .B1(n4481), .B2(n568), .ZN(n4696)
         );
  NAND2_X1 U3529 ( .A1(n4698), .A2(n4699), .ZN(n4691) );
  AOI22_X1 U3530 ( .A1(n5596), .A2(n696), .B1(n5591), .B2(n664), .ZN(n4699) );
  AOI22_X1 U3531 ( .A1(n5590), .A2(n728), .B1(n5587), .B2(n600), .ZN(n4698) );
  NAND2_X1 U3532 ( .A1(n4700), .A2(n4701), .ZN(n4690) );
  AOI22_X1 U3533 ( .A1(n5584), .A2(n504), .B1(n5581), .B2(n376), .ZN(n4701) );
  AOI22_X1 U3534 ( .A1(n5578), .A2(n536), .B1(n5573), .B2(n344), .ZN(n4700) );
  NAND2_X1 U3535 ( .A1(n4702), .A2(n4703), .ZN(n3188) );
  NOR4_X1 U3536 ( .A1(n4704), .A2(n4705), .A3(n4706), .A4(n4707), .ZN(n4703)
         );
  OAI21_X1 U3537 ( .B1(n1432), .B2(n5668), .A(n4708), .ZN(n4707) );
  NAND2_X1 U3538 ( .A1(n4444), .A2(n6461), .ZN(n4708) );
  OAI21_X1 U3539 ( .B1(n6085), .B2(n5662), .A(n4709), .ZN(n4706) );
  AOI22_X1 U3540 ( .A1(n5659), .A2(n6397), .B1(n5656), .B2(n6429), .ZN(n4709)
         );
  NAND2_X1 U3541 ( .A1(n4710), .A2(n4711), .ZN(n4705) );
  AOI22_X1 U3542 ( .A1(n5653), .A2(n2821), .B1(n5650), .B2(n6525), .ZN(n4711)
         );
  AOI22_X1 U3543 ( .A1(n5645), .A2(n6365), .B1(n5644), .B2(n6565), .ZN(n4710)
         );
  AOI22_X1 U3545 ( .A1(n5641), .A2(n2355), .B1(n5638), .B2(n6312), .ZN(n4715)
         );
  AOI22_X1 U3546 ( .A1(n4461), .A2(n6149), .B1(n5632), .B2(n6597), .ZN(n4714)
         );
  AOI22_X1 U3547 ( .A1(n5629), .A2(n2240), .B1(n5626), .B2(n6248), .ZN(n4713)
         );
  AOI22_X1 U3548 ( .A1(n5623), .A2(n631), .B1(n5620), .B2(n471), .ZN(n4712) );
  NOR4_X1 U3549 ( .A1(n4716), .A2(n4717), .A3(n4718), .A4(n4719), .ZN(n4702)
         );
  NAND2_X1 U3550 ( .A1(n4720), .A2(n4721), .ZN(n4719) );
  AOI22_X1 U3551 ( .A1(n5617), .A2(n407), .B1(n5614), .B2(n6181), .ZN(n4721)
         );
  AOI22_X1 U3552 ( .A1(n5611), .A2(n6280), .B1(n5457), .B2(OUT2[22]), .ZN(
        n4720) );
  NAND2_X1 U3553 ( .A1(n4722), .A2(n4723), .ZN(n4718) );
  AOI22_X1 U3554 ( .A1(n5608), .A2(n439), .B1(n5605), .B2(n6117), .ZN(n4723)
         );
  AOI22_X1 U3555 ( .A1(n5602), .A2(n6213), .B1(n4481), .B2(n567), .ZN(n4722)
         );
  NAND2_X1 U3556 ( .A1(n4724), .A2(n4725), .ZN(n4717) );
  AOI22_X1 U3557 ( .A1(n5596), .A2(n695), .B1(n5591), .B2(n663), .ZN(n4725) );
  AOI22_X1 U3558 ( .A1(n5590), .A2(n727), .B1(n5587), .B2(n599), .ZN(n4724) );
  NAND2_X1 U3559 ( .A1(n4726), .A2(n4727), .ZN(n4716) );
  AOI22_X1 U3560 ( .A1(n5584), .A2(n503), .B1(n5581), .B2(n375), .ZN(n4727) );
  AOI22_X1 U3561 ( .A1(n5578), .A2(n535), .B1(n5573), .B2(n343), .ZN(n4726) );
  NAND2_X1 U3562 ( .A1(n4728), .A2(n4729), .ZN(n3187) );
  NOR4_X1 U3563 ( .A1(n4730), .A2(n4731), .A3(n4732), .A4(n4733), .ZN(n4729)
         );
  OAI21_X1 U3564 ( .B1(n1433), .B2(n4442), .A(n4734), .ZN(n4733) );
  NAND2_X1 U3565 ( .A1(n5664), .A2(n6462), .ZN(n4734) );
  OAI21_X1 U3566 ( .B1(n6086), .B2(n4445), .A(n4735), .ZN(n4732) );
  AOI22_X1 U3567 ( .A1(n5659), .A2(n6398), .B1(n5656), .B2(n6430), .ZN(n4735)
         );
  NAND2_X1 U3568 ( .A1(n4736), .A2(n4737), .ZN(n4731) );
  AOI22_X1 U3569 ( .A1(n4451), .A2(n2820), .B1(n5650), .B2(n6526), .ZN(n4737)
         );
  AOI22_X1 U3570 ( .A1(n5645), .A2(n6366), .B1(n5644), .B2(n6566), .ZN(n4736)
         );
  AOI22_X1 U3572 ( .A1(n5641), .A2(n2352), .B1(n5638), .B2(n6313), .ZN(n4741)
         );
  AOI22_X1 U3573 ( .A1(n5634), .A2(n6150), .B1(n5632), .B2(n6598), .ZN(n4740)
         );
  AOI22_X1 U3574 ( .A1(n5629), .A2(n2235), .B1(n5626), .B2(n6249), .ZN(n4739)
         );
  AOI22_X1 U3575 ( .A1(n5623), .A2(n630), .B1(n5620), .B2(n470), .ZN(n4738) );
  NOR4_X1 U3576 ( .A1(n4742), .A2(n4743), .A3(n4744), .A4(n4745), .ZN(n4728)
         );
  NAND2_X1 U3577 ( .A1(n4746), .A2(n4747), .ZN(n4745) );
  AOI22_X1 U3578 ( .A1(n5617), .A2(n406), .B1(n5614), .B2(n6182), .ZN(n4747)
         );
  AOI22_X1 U3579 ( .A1(n5611), .A2(n6281), .B1(n5457), .B2(OUT2[21]), .ZN(
        n4746) );
  NAND2_X1 U3580 ( .A1(n4748), .A2(n4749), .ZN(n4744) );
  AOI22_X1 U3581 ( .A1(n5608), .A2(n438), .B1(n5605), .B2(n6118), .ZN(n4749)
         );
  AOI22_X1 U3582 ( .A1(n5602), .A2(n6214), .B1(n5598), .B2(n566), .ZN(n4748)
         );
  NAND2_X1 U3583 ( .A1(n4750), .A2(n4751), .ZN(n4743) );
  AOI22_X1 U3584 ( .A1(n5596), .A2(n694), .B1(n4485), .B2(n662), .ZN(n4751) );
  AOI22_X1 U3585 ( .A1(n5590), .A2(n726), .B1(n5587), .B2(n598), .ZN(n4750) );
  NAND2_X1 U3586 ( .A1(n4752), .A2(n4753), .ZN(n4742) );
  AOI22_X1 U3587 ( .A1(n5584), .A2(n502), .B1(n5581), .B2(n374), .ZN(n4753) );
  AOI22_X1 U3588 ( .A1(n5578), .A2(n534), .B1(n4493), .B2(n342), .ZN(n4752) );
  NAND2_X1 U3589 ( .A1(n4754), .A2(n4755), .ZN(n3186) );
  NOR4_X1 U3590 ( .A1(n4756), .A2(n4757), .A3(n4758), .A4(n4759), .ZN(n4755)
         );
  OAI21_X1 U3591 ( .B1(n1434), .B2(n4442), .A(n4760), .ZN(n4759) );
  NAND2_X1 U3592 ( .A1(n5664), .A2(n6463), .ZN(n4760) );
  OAI21_X1 U3593 ( .B1(n6087), .B2(n4445), .A(n4761), .ZN(n4758) );
  AOI22_X1 U3594 ( .A1(n5659), .A2(n6399), .B1(n5656), .B2(n6431), .ZN(n4761)
         );
  NAND2_X1 U3595 ( .A1(n4762), .A2(n4763), .ZN(n4757) );
  AOI22_X1 U3596 ( .A1(n5653), .A2(n2819), .B1(n5650), .B2(n6527), .ZN(n4763)
         );
  AOI22_X1 U3597 ( .A1(n4453), .A2(n6367), .B1(n5644), .B2(n6567), .ZN(n4762)
         );
  AOI22_X1 U3599 ( .A1(n5641), .A2(n6335), .B1(n5638), .B2(n6314), .ZN(n4767)
         );
  AOI22_X1 U3600 ( .A1(n5634), .A2(n6151), .B1(n5632), .B2(n6599), .ZN(n4766)
         );
  AOI22_X1 U3601 ( .A1(n5629), .A2(n2230), .B1(n5626), .B2(n6250), .ZN(n4765)
         );
  AOI22_X1 U3602 ( .A1(n5623), .A2(n629), .B1(n5620), .B2(n469), .ZN(n4764) );
  NOR4_X1 U3603 ( .A1(n4768), .A2(n4769), .A3(n4770), .A4(n4771), .ZN(n4754)
         );
  NAND2_X1 U3604 ( .A1(n4772), .A2(n4773), .ZN(n4771) );
  AOI22_X1 U3605 ( .A1(n5617), .A2(n405), .B1(n5614), .B2(n6183), .ZN(n4773)
         );
  AOI22_X1 U3606 ( .A1(n5611), .A2(n6282), .B1(n5457), .B2(OUT2[20]), .ZN(
        n4772) );
  NAND2_X1 U3607 ( .A1(n4774), .A2(n4775), .ZN(n4770) );
  AOI22_X1 U3608 ( .A1(n5608), .A2(n437), .B1(n5605), .B2(n6119), .ZN(n4775)
         );
  AOI22_X1 U3609 ( .A1(n5602), .A2(n6215), .B1(n5598), .B2(n565), .ZN(n4774)
         );
  NAND2_X1 U3610 ( .A1(n4776), .A2(n4777), .ZN(n4769) );
  AOI22_X1 U3611 ( .A1(n5596), .A2(n693), .B1(n4485), .B2(n661), .ZN(n4777) );
  AOI22_X1 U3612 ( .A1(n5590), .A2(n725), .B1(n5587), .B2(n597), .ZN(n4776) );
  NAND2_X1 U3613 ( .A1(n4778), .A2(n4779), .ZN(n4768) );
  AOI22_X1 U3614 ( .A1(n5584), .A2(n501), .B1(n5581), .B2(n373), .ZN(n4779) );
  AOI22_X1 U3615 ( .A1(n5578), .A2(n533), .B1(n4493), .B2(n341), .ZN(n4778) );
  NAND2_X1 U3616 ( .A1(n4780), .A2(n4781), .ZN(n3185) );
  NOR4_X1 U3617 ( .A1(n4782), .A2(n4783), .A3(n4784), .A4(n4785), .ZN(n4781)
         );
  OAI21_X1 U3618 ( .B1(n1435), .B2(n4442), .A(n4786), .ZN(n4785) );
  NAND2_X1 U3619 ( .A1(n5664), .A2(n6464), .ZN(n4786) );
  OAI21_X1 U3620 ( .B1(n6088), .B2(n4445), .A(n4787), .ZN(n4784) );
  AOI22_X1 U3621 ( .A1(n5659), .A2(n6400), .B1(n5656), .B2(n6432), .ZN(n4787)
         );
  NAND2_X1 U3622 ( .A1(n4788), .A2(n4789), .ZN(n4783) );
  AOI22_X1 U3623 ( .A1(n5653), .A2(n2818), .B1(n5650), .B2(n6528), .ZN(n4789)
         );
  AOI22_X1 U3624 ( .A1(n4453), .A2(n6368), .B1(n5644), .B2(n6568), .ZN(n4788)
         );
  AOI22_X1 U3626 ( .A1(n5641), .A2(n6336), .B1(n5638), .B2(n6315), .ZN(n4793)
         );
  AOI22_X1 U3627 ( .A1(n5634), .A2(n6152), .B1(n5632), .B2(n6600), .ZN(n4792)
         );
  AOI22_X1 U3628 ( .A1(n5629), .A2(n2225), .B1(n5626), .B2(n6251), .ZN(n4791)
         );
  AOI22_X1 U3629 ( .A1(n5623), .A2(n628), .B1(n5620), .B2(n468), .ZN(n4790) );
  NOR4_X1 U3630 ( .A1(n4794), .A2(n4795), .A3(n4796), .A4(n4797), .ZN(n4780)
         );
  NAND2_X1 U3631 ( .A1(n4798), .A2(n4799), .ZN(n4797) );
  AOI22_X1 U3632 ( .A1(n5617), .A2(n404), .B1(n5614), .B2(n6184), .ZN(n4799)
         );
  AOI22_X1 U3633 ( .A1(n5611), .A2(n6283), .B1(n5458), .B2(OUT2[19]), .ZN(
        n4798) );
  NAND2_X1 U3634 ( .A1(n4800), .A2(n4801), .ZN(n4796) );
  AOI22_X1 U3635 ( .A1(n5608), .A2(n436), .B1(n5605), .B2(n6120), .ZN(n4801)
         );
  AOI22_X1 U3636 ( .A1(n5602), .A2(n6216), .B1(n5598), .B2(n564), .ZN(n4800)
         );
  NAND2_X1 U3637 ( .A1(n4802), .A2(n4803), .ZN(n4795) );
  AOI22_X1 U3638 ( .A1(n5596), .A2(n692), .B1(n4485), .B2(n660), .ZN(n4803) );
  AOI22_X1 U3639 ( .A1(n5590), .A2(n724), .B1(n5587), .B2(n596), .ZN(n4802) );
  NAND2_X1 U3640 ( .A1(n4804), .A2(n4805), .ZN(n4794) );
  AOI22_X1 U3641 ( .A1(n5584), .A2(n500), .B1(n5581), .B2(n372), .ZN(n4805) );
  AOI22_X1 U3642 ( .A1(n5578), .A2(n532), .B1(n4493), .B2(n340), .ZN(n4804) );
  NAND2_X1 U3643 ( .A1(n4806), .A2(n4807), .ZN(n3184) );
  NOR4_X1 U3644 ( .A1(n4808), .A2(n4809), .A3(n4810), .A4(n4811), .ZN(n4807)
         );
  OAI21_X1 U3645 ( .B1(n1436), .B2(n4442), .A(n4812), .ZN(n4811) );
  NAND2_X1 U3646 ( .A1(n5664), .A2(n6465), .ZN(n4812) );
  OAI21_X1 U3647 ( .B1(n6089), .B2(n4445), .A(n4813), .ZN(n4810) );
  AOI22_X1 U3648 ( .A1(n5659), .A2(n6401), .B1(n5656), .B2(n6433), .ZN(n4813)
         );
  NAND2_X1 U3649 ( .A1(n4814), .A2(n4815), .ZN(n4809) );
  AOI22_X1 U3650 ( .A1(n5653), .A2(n2817), .B1(n5650), .B2(n6529), .ZN(n4815)
         );
  AOI22_X1 U3651 ( .A1(n4453), .A2(n6369), .B1(n5644), .B2(n6569), .ZN(n4814)
         );
  AOI22_X1 U3653 ( .A1(n5641), .A2(n6337), .B1(n5638), .B2(n6316), .ZN(n4819)
         );
  AOI22_X1 U3654 ( .A1(n5634), .A2(n6153), .B1(n5632), .B2(n6601), .ZN(n4818)
         );
  AOI22_X1 U3655 ( .A1(n5629), .A2(n2220), .B1(n5626), .B2(n6252), .ZN(n4817)
         );
  AOI22_X1 U3656 ( .A1(n5623), .A2(n627), .B1(n5620), .B2(n467), .ZN(n4816) );
  NOR4_X1 U3657 ( .A1(n4820), .A2(n4821), .A3(n4822), .A4(n4823), .ZN(n4806)
         );
  NAND2_X1 U3658 ( .A1(n4824), .A2(n4825), .ZN(n4823) );
  AOI22_X1 U3659 ( .A1(n5617), .A2(n403), .B1(n5614), .B2(n6185), .ZN(n4825)
         );
  AOI22_X1 U3660 ( .A1(n5611), .A2(n6284), .B1(n5457), .B2(OUT2[18]), .ZN(
        n4824) );
  NAND2_X1 U3661 ( .A1(n4826), .A2(n4827), .ZN(n4822) );
  AOI22_X1 U3662 ( .A1(n5608), .A2(n435), .B1(n5605), .B2(n6121), .ZN(n4827)
         );
  AOI22_X1 U3663 ( .A1(n5602), .A2(n6217), .B1(n5598), .B2(n563), .ZN(n4826)
         );
  NAND2_X1 U3664 ( .A1(n4828), .A2(n4829), .ZN(n4821) );
  AOI22_X1 U3665 ( .A1(n5596), .A2(n691), .B1(n4485), .B2(n659), .ZN(n4829) );
  AOI22_X1 U3666 ( .A1(n5590), .A2(n723), .B1(n5587), .B2(n595), .ZN(n4828) );
  NAND2_X1 U3667 ( .A1(n4830), .A2(n4831), .ZN(n4820) );
  AOI22_X1 U3668 ( .A1(n5584), .A2(n499), .B1(n5581), .B2(n371), .ZN(n4831) );
  AOI22_X1 U3669 ( .A1(n5578), .A2(n531), .B1(n4493), .B2(n339), .ZN(n4830) );
  NAND2_X1 U3670 ( .A1(n4832), .A2(n4833), .ZN(n3183) );
  NOR4_X1 U3671 ( .A1(n4834), .A2(n4835), .A3(n4836), .A4(n4837), .ZN(n4833)
         );
  OAI21_X1 U3672 ( .B1(n1437), .B2(n4442), .A(n4838), .ZN(n4837) );
  NAND2_X1 U3673 ( .A1(n5664), .A2(n6466), .ZN(n4838) );
  OAI21_X1 U3674 ( .B1(n6090), .B2(n4445), .A(n4839), .ZN(n4836) );
  AOI22_X1 U3675 ( .A1(n5659), .A2(n6402), .B1(n5656), .B2(n6434), .ZN(n4839)
         );
  NAND2_X1 U3676 ( .A1(n4840), .A2(n4841), .ZN(n4835) );
  AOI22_X1 U3677 ( .A1(n5653), .A2(n2816), .B1(n5650), .B2(n6530), .ZN(n4841)
         );
  AOI22_X1 U3678 ( .A1(n4453), .A2(n6370), .B1(n5644), .B2(n6570), .ZN(n4840)
         );
  AOI22_X1 U3680 ( .A1(n5641), .A2(n6338), .B1(n5638), .B2(n6317), .ZN(n4845)
         );
  AOI22_X1 U3681 ( .A1(n5634), .A2(n6154), .B1(n5632), .B2(n6602), .ZN(n4844)
         );
  AOI22_X1 U3682 ( .A1(n5629), .A2(n2215), .B1(n5626), .B2(n6253), .ZN(n4843)
         );
  AOI22_X1 U3683 ( .A1(n5623), .A2(n626), .B1(n5620), .B2(n466), .ZN(n4842) );
  NOR4_X1 U3684 ( .A1(n4846), .A2(n4847), .A3(n4848), .A4(n4849), .ZN(n4832)
         );
  NAND2_X1 U3685 ( .A1(n4850), .A2(n4851), .ZN(n4849) );
  AOI22_X1 U3686 ( .A1(n5617), .A2(n402), .B1(n5614), .B2(n6186), .ZN(n4851)
         );
  AOI22_X1 U3687 ( .A1(n5611), .A2(n6285), .B1(n5457), .B2(OUT2[17]), .ZN(
        n4850) );
  NAND2_X1 U3688 ( .A1(n4852), .A2(n4853), .ZN(n4848) );
  AOI22_X1 U3689 ( .A1(n5608), .A2(n434), .B1(n5605), .B2(n6122), .ZN(n4853)
         );
  AOI22_X1 U3690 ( .A1(n5602), .A2(n6218), .B1(n5598), .B2(n562), .ZN(n4852)
         );
  NAND2_X1 U3691 ( .A1(n4854), .A2(n4855), .ZN(n4847) );
  AOI22_X1 U3692 ( .A1(n5596), .A2(n690), .B1(n4485), .B2(n658), .ZN(n4855) );
  AOI22_X1 U3693 ( .A1(n5590), .A2(n722), .B1(n5587), .B2(n594), .ZN(n4854) );
  NAND2_X1 U3694 ( .A1(n4856), .A2(n4857), .ZN(n4846) );
  AOI22_X1 U3695 ( .A1(n5584), .A2(n498), .B1(n5581), .B2(n370), .ZN(n4857) );
  AOI22_X1 U3696 ( .A1(n5578), .A2(n530), .B1(n4493), .B2(n338), .ZN(n4856) );
  NAND2_X1 U3697 ( .A1(n4858), .A2(n4859), .ZN(n3182) );
  NOR4_X1 U3698 ( .A1(n4860), .A2(n4861), .A3(n4862), .A4(n4863), .ZN(n4859)
         );
  OAI21_X1 U3699 ( .B1(n1438), .B2(n4442), .A(n4864), .ZN(n4863) );
  NAND2_X1 U3700 ( .A1(n5664), .A2(n6467), .ZN(n4864) );
  OAI21_X1 U3701 ( .B1(n6091), .B2(n4445), .A(n4865), .ZN(n4862) );
  AOI22_X1 U3702 ( .A1(n5659), .A2(n6403), .B1(n5656), .B2(n6435), .ZN(n4865)
         );
  NAND2_X1 U3703 ( .A1(n4866), .A2(n4867), .ZN(n4861) );
  AOI22_X1 U3704 ( .A1(n5653), .A2(n2815), .B1(n5650), .B2(n6531), .ZN(n4867)
         );
  AOI22_X1 U3705 ( .A1(n4453), .A2(n6371), .B1(n5644), .B2(n6571), .ZN(n4866)
         );
  AOI22_X1 U3707 ( .A1(n5641), .A2(n6339), .B1(n5638), .B2(n6318), .ZN(n4871)
         );
  AOI22_X1 U3708 ( .A1(n5634), .A2(n6155), .B1(n5632), .B2(n6603), .ZN(n4870)
         );
  AOI22_X1 U3709 ( .A1(n5629), .A2(n2210), .B1(n5626), .B2(n6254), .ZN(n4869)
         );
  AOI22_X1 U3710 ( .A1(n5623), .A2(n625), .B1(n5620), .B2(n465), .ZN(n4868) );
  NOR4_X1 U3711 ( .A1(n4872), .A2(n4873), .A3(n4874), .A4(n4875), .ZN(n4858)
         );
  NAND2_X1 U3712 ( .A1(n4876), .A2(n4877), .ZN(n4875) );
  AOI22_X1 U3713 ( .A1(n5617), .A2(n401), .B1(n5614), .B2(n6187), .ZN(n4877)
         );
  AOI22_X1 U3714 ( .A1(n5611), .A2(n6286), .B1(n5457), .B2(OUT2[16]), .ZN(
        n4876) );
  NAND2_X1 U3715 ( .A1(n4878), .A2(n4879), .ZN(n4874) );
  AOI22_X1 U3716 ( .A1(n5608), .A2(n433), .B1(n5605), .B2(n6123), .ZN(n4879)
         );
  AOI22_X1 U3717 ( .A1(n5602), .A2(n6219), .B1(n5598), .B2(n561), .ZN(n4878)
         );
  NAND2_X1 U3718 ( .A1(n4880), .A2(n4881), .ZN(n4873) );
  AOI22_X1 U3719 ( .A1(n5596), .A2(n689), .B1(n4485), .B2(n657), .ZN(n4881) );
  AOI22_X1 U3720 ( .A1(n5590), .A2(n721), .B1(n5587), .B2(n593), .ZN(n4880) );
  NAND2_X1 U3721 ( .A1(n4882), .A2(n4883), .ZN(n4872) );
  AOI22_X1 U3722 ( .A1(n5584), .A2(n497), .B1(n5581), .B2(n369), .ZN(n4883) );
  AOI22_X1 U3723 ( .A1(n5578), .A2(n529), .B1(n4493), .B2(n337), .ZN(n4882) );
  NAND2_X1 U3724 ( .A1(n4884), .A2(n4885), .ZN(n3181) );
  NOR4_X1 U3725 ( .A1(n4886), .A2(n4887), .A3(n4888), .A4(n4889), .ZN(n4885)
         );
  OAI21_X1 U3726 ( .B1(n1439), .B2(n4442), .A(n4890), .ZN(n4889) );
  NAND2_X1 U3727 ( .A1(n5664), .A2(n6468), .ZN(n4890) );
  OAI21_X1 U3728 ( .B1(n5507), .B2(n4445), .A(n4891), .ZN(n4888) );
  AOI22_X1 U3729 ( .A1(n5659), .A2(n6404), .B1(n5656), .B2(n6436), .ZN(n4891)
         );
  NAND2_X1 U3730 ( .A1(n4892), .A2(n4893), .ZN(n4887) );
  AOI22_X1 U3731 ( .A1(n5653), .A2(n2814), .B1(n5650), .B2(n6532), .ZN(n4893)
         );
  AOI22_X1 U3732 ( .A1(n4453), .A2(n6372), .B1(n5644), .B2(n6572), .ZN(n4892)
         );
  AOI22_X1 U3734 ( .A1(n5641), .A2(n6340), .B1(n5638), .B2(n6319), .ZN(n4897)
         );
  AOI22_X1 U3735 ( .A1(n5634), .A2(n6156), .B1(n5632), .B2(n6604), .ZN(n4896)
         );
  AOI22_X1 U3736 ( .A1(n5629), .A2(n2205), .B1(n5626), .B2(n6255), .ZN(n4895)
         );
  AOI22_X1 U3737 ( .A1(n5623), .A2(n624), .B1(n5620), .B2(n464), .ZN(n4894) );
  NOR4_X1 U3738 ( .A1(n4898), .A2(n4899), .A3(n4900), .A4(n4901), .ZN(n4884)
         );
  NAND2_X1 U3739 ( .A1(n4902), .A2(n4903), .ZN(n4901) );
  AOI22_X1 U3740 ( .A1(n5617), .A2(n400), .B1(n5614), .B2(n6188), .ZN(n4903)
         );
  AOI22_X1 U3741 ( .A1(n5611), .A2(n6287), .B1(n5458), .B2(OUT2[15]), .ZN(
        n4902) );
  NAND2_X1 U3742 ( .A1(n4904), .A2(n4905), .ZN(n4900) );
  AOI22_X1 U3743 ( .A1(n5608), .A2(n432), .B1(n5605), .B2(n6124), .ZN(n4905)
         );
  AOI22_X1 U3744 ( .A1(n5602), .A2(n6220), .B1(n5598), .B2(n560), .ZN(n4904)
         );
  NAND2_X1 U3745 ( .A1(n4906), .A2(n4907), .ZN(n4899) );
  AOI22_X1 U3746 ( .A1(n5596), .A2(n688), .B1(n4485), .B2(n656), .ZN(n4907) );
  AOI22_X1 U3747 ( .A1(n5590), .A2(n720), .B1(n5587), .B2(n592), .ZN(n4906) );
  NAND2_X1 U3748 ( .A1(n4908), .A2(n4909), .ZN(n4898) );
  AOI22_X1 U3749 ( .A1(n5584), .A2(n496), .B1(n5581), .B2(n368), .ZN(n4909) );
  AOI22_X1 U3750 ( .A1(n5578), .A2(n528), .B1(n4493), .B2(n336), .ZN(n4908) );
  NAND2_X1 U3751 ( .A1(n4910), .A2(n4911), .ZN(n3180) );
  NOR4_X1 U3752 ( .A1(n4912), .A2(n4913), .A3(n4914), .A4(n4915), .ZN(n4911)
         );
  OAI21_X1 U3753 ( .B1(n1440), .B2(n4442), .A(n4916), .ZN(n4915) );
  NAND2_X1 U3754 ( .A1(n5664), .A2(n6469), .ZN(n4916) );
  OAI21_X1 U3755 ( .B1(n6093), .B2(n4445), .A(n4917), .ZN(n4914) );
  AOI22_X1 U3756 ( .A1(n5659), .A2(n6405), .B1(n5656), .B2(n6437), .ZN(n4917)
         );
  NAND2_X1 U3757 ( .A1(n4918), .A2(n4919), .ZN(n4913) );
  AOI22_X1 U3758 ( .A1(n5653), .A2(n2813), .B1(n5650), .B2(n6533), .ZN(n4919)
         );
  AOI22_X1 U3759 ( .A1(n4453), .A2(n6373), .B1(n5644), .B2(n6573), .ZN(n4918)
         );
  AOI22_X1 U3761 ( .A1(n5641), .A2(n6341), .B1(n5638), .B2(n6320), .ZN(n4923)
         );
  AOI22_X1 U3762 ( .A1(n5634), .A2(n6157), .B1(n5632), .B2(n6605), .ZN(n4922)
         );
  AOI22_X1 U3763 ( .A1(n5629), .A2(n2200), .B1(n5626), .B2(n6256), .ZN(n4921)
         );
  AOI22_X1 U3764 ( .A1(n5623), .A2(n623), .B1(n5620), .B2(n463), .ZN(n4920) );
  NOR4_X1 U3765 ( .A1(n4924), .A2(n4925), .A3(n4926), .A4(n4927), .ZN(n4910)
         );
  NAND2_X1 U3766 ( .A1(n4928), .A2(n4929), .ZN(n4927) );
  AOI22_X1 U3767 ( .A1(n5617), .A2(n399), .B1(n5614), .B2(n6189), .ZN(n4929)
         );
  AOI22_X1 U3768 ( .A1(n5611), .A2(n6288), .B1(n5457), .B2(OUT2[14]), .ZN(
        n4928) );
  NAND2_X1 U3769 ( .A1(n4930), .A2(n4931), .ZN(n4926) );
  AOI22_X1 U3770 ( .A1(n5608), .A2(n431), .B1(n5605), .B2(n6125), .ZN(n4931)
         );
  AOI22_X1 U3771 ( .A1(n5602), .A2(n6221), .B1(n5598), .B2(n559), .ZN(n4930)
         );
  NAND2_X1 U3772 ( .A1(n4932), .A2(n4933), .ZN(n4925) );
  AOI22_X1 U3773 ( .A1(n5596), .A2(n687), .B1(n4485), .B2(n655), .ZN(n4933) );
  AOI22_X1 U3774 ( .A1(n5590), .A2(n719), .B1(n5587), .B2(n591), .ZN(n4932) );
  NAND2_X1 U3775 ( .A1(n4934), .A2(n4935), .ZN(n4924) );
  AOI22_X1 U3776 ( .A1(n5584), .A2(n495), .B1(n5581), .B2(n367), .ZN(n4935) );
  AOI22_X1 U3777 ( .A1(n5578), .A2(n527), .B1(n4493), .B2(n335), .ZN(n4934) );
  NAND2_X1 U3778 ( .A1(n4936), .A2(n4937), .ZN(n3179) );
  NOR4_X1 U3779 ( .A1(n4938), .A2(n4939), .A3(n4940), .A4(n4941), .ZN(n4937)
         );
  OAI21_X1 U3780 ( .B1(n1441), .B2(n4442), .A(n4942), .ZN(n4941) );
  NAND2_X1 U3781 ( .A1(n5664), .A2(n6470), .ZN(n4942) );
  OAI21_X1 U3782 ( .B1(n6094), .B2(n4445), .A(n4943), .ZN(n4940) );
  AOI22_X1 U3783 ( .A1(n5659), .A2(n6406), .B1(n5656), .B2(n6438), .ZN(n4943)
         );
  NAND2_X1 U3784 ( .A1(n4944), .A2(n4945), .ZN(n4939) );
  AOI22_X1 U3785 ( .A1(n5653), .A2(n2812), .B1(n5650), .B2(n6534), .ZN(n4945)
         );
  AOI22_X1 U3786 ( .A1(n4453), .A2(n6374), .B1(n5644), .B2(n6574), .ZN(n4944)
         );
  AOI22_X1 U3788 ( .A1(n5641), .A2(n6342), .B1(n5638), .B2(n6321), .ZN(n4949)
         );
  AOI22_X1 U3789 ( .A1(n5634), .A2(n6158), .B1(n5632), .B2(n6606), .ZN(n4948)
         );
  AOI22_X1 U3790 ( .A1(n5629), .A2(n2195), .B1(n5626), .B2(n6257), .ZN(n4947)
         );
  AOI22_X1 U3791 ( .A1(n5623), .A2(n622), .B1(n5620), .B2(n462), .ZN(n4946) );
  NOR4_X1 U3792 ( .A1(n4950), .A2(n4951), .A3(n4952), .A4(n4953), .ZN(n4936)
         );
  NAND2_X1 U3793 ( .A1(n4954), .A2(n4955), .ZN(n4953) );
  AOI22_X1 U3794 ( .A1(n4473), .A2(n398), .B1(n5614), .B2(n6190), .ZN(n4955)
         );
  AOI22_X1 U3795 ( .A1(n4475), .A2(n6289), .B1(n5458), .B2(OUT2[13]), .ZN(
        n4954) );
  NAND2_X1 U3796 ( .A1(n4956), .A2(n4957), .ZN(n4952) );
  AOI22_X1 U3797 ( .A1(n4478), .A2(n430), .B1(n5605), .B2(n6126), .ZN(n4957)
         );
  AOI22_X1 U3798 ( .A1(n5602), .A2(n6222), .B1(n5598), .B2(n558), .ZN(n4956)
         );
  NAND2_X1 U3799 ( .A1(n4958), .A2(n4959), .ZN(n4951) );
  AOI22_X1 U3800 ( .A1(n4484), .A2(n686), .B1(n4485), .B2(n654), .ZN(n4959) );
  AOI22_X1 U3801 ( .A1(n5590), .A2(n718), .B1(n5587), .B2(n590), .ZN(n4958) );
  NAND2_X1 U3802 ( .A1(n4960), .A2(n4961), .ZN(n4950) );
  AOI22_X1 U3803 ( .A1(n4490), .A2(n494), .B1(n5581), .B2(n366), .ZN(n4961) );
  AOI22_X1 U3804 ( .A1(n5578), .A2(n526), .B1(n4493), .B2(n334), .ZN(n4960) );
  NAND2_X1 U3805 ( .A1(n4962), .A2(n4963), .ZN(n3178) );
  NOR4_X1 U3806 ( .A1(n4964), .A2(n4965), .A3(n4966), .A4(n4967), .ZN(n4963)
         );
  OAI21_X1 U3807 ( .B1(n1442), .B2(n4442), .A(n4968), .ZN(n4967) );
  NAND2_X1 U3808 ( .A1(n5664), .A2(n6471), .ZN(n4968) );
  OAI21_X1 U3809 ( .B1(n6095), .B2(n4445), .A(n4969), .ZN(n4966) );
  AOI22_X1 U3810 ( .A1(n4447), .A2(n6407), .B1(n5656), .B2(n6439), .ZN(n4969)
         );
  NAND2_X1 U3811 ( .A1(n4970), .A2(n4971), .ZN(n4965) );
  AOI22_X1 U3812 ( .A1(n5653), .A2(n2811), .B1(n5650), .B2(n6535), .ZN(n4971)
         );
  AOI22_X1 U3813 ( .A1(n4453), .A2(n6375), .B1(n5644), .B2(n6575), .ZN(n4970)
         );
  AOI22_X1 U3815 ( .A1(n4459), .A2(n6343), .B1(n5638), .B2(n6322), .ZN(n4975)
         );
  AOI22_X1 U3816 ( .A1(n5634), .A2(n6159), .B1(n5632), .B2(n6607), .ZN(n4974)
         );
  AOI22_X1 U3817 ( .A1(n4463), .A2(n2190), .B1(n5626), .B2(n6258), .ZN(n4973)
         );
  AOI22_X1 U3818 ( .A1(n4465), .A2(n621), .B1(n5620), .B2(n461), .ZN(n4972) );
  NOR4_X1 U3819 ( .A1(n4976), .A2(n4977), .A3(n4978), .A4(n4979), .ZN(n4962)
         );
  NAND2_X1 U3820 ( .A1(n4980), .A2(n4981), .ZN(n4979) );
  AOI22_X1 U3821 ( .A1(n5617), .A2(n397), .B1(n5614), .B2(n6191), .ZN(n4981)
         );
  AOI22_X1 U3822 ( .A1(n5611), .A2(n6290), .B1(n5457), .B2(OUT2[12]), .ZN(
        n4980) );
  NAND2_X1 U3823 ( .A1(n4982), .A2(n4983), .ZN(n4978) );
  AOI22_X1 U3824 ( .A1(n5608), .A2(n429), .B1(n5605), .B2(n6127), .ZN(n4983)
         );
  AOI22_X1 U3825 ( .A1(n4480), .A2(n6223), .B1(n5598), .B2(n557), .ZN(n4982)
         );
  NAND2_X1 U3826 ( .A1(n4984), .A2(n4985), .ZN(n4977) );
  AOI22_X1 U3827 ( .A1(n5596), .A2(n685), .B1(n4485), .B2(n653), .ZN(n4985) );
  AOI22_X1 U3828 ( .A1(n4486), .A2(n717), .B1(n5587), .B2(n589), .ZN(n4984) );
  NAND2_X1 U3829 ( .A1(n4986), .A2(n4987), .ZN(n4976) );
  AOI22_X1 U3830 ( .A1(n5584), .A2(n493), .B1(n5581), .B2(n365), .ZN(n4987) );
  AOI22_X1 U3831 ( .A1(n4492), .A2(n525), .B1(n4493), .B2(n333), .ZN(n4986) );
  NAND2_X1 U3832 ( .A1(n4988), .A2(n4989), .ZN(n3177) );
  NOR4_X1 U3833 ( .A1(n4990), .A2(n4991), .A3(n4992), .A4(n4993), .ZN(n4989)
         );
  OAI21_X1 U3834 ( .B1(n1443), .B2(n4442), .A(n4994), .ZN(n4993) );
  NAND2_X1 U3835 ( .A1(n5664), .A2(n6472), .ZN(n4994) );
  OAI21_X1 U3836 ( .B1(n6096), .B2(n4445), .A(n4995), .ZN(n4992) );
  AOI22_X1 U3837 ( .A1(n5659), .A2(n6408), .B1(n5656), .B2(n6440), .ZN(n4995)
         );
  NAND2_X1 U3838 ( .A1(n4996), .A2(n4997), .ZN(n4991) );
  AOI22_X1 U3839 ( .A1(n5653), .A2(n2810), .B1(n5650), .B2(n6536), .ZN(n4997)
         );
  AOI22_X1 U3840 ( .A1(n5645), .A2(n6376), .B1(n5644), .B2(n6576), .ZN(n4996)
         );
  AOI22_X1 U3842 ( .A1(n5641), .A2(n6344), .B1(n5638), .B2(n6323), .ZN(n5001)
         );
  AOI22_X1 U3843 ( .A1(n5634), .A2(n6160), .B1(n5632), .B2(n6608), .ZN(n5000)
         );
  AOI22_X1 U3844 ( .A1(n5629), .A2(n2185), .B1(n5626), .B2(n6259), .ZN(n4999)
         );
  AOI22_X1 U3845 ( .A1(n5623), .A2(n620), .B1(n5620), .B2(n460), .ZN(n4998) );
  NOR4_X1 U3846 ( .A1(n5002), .A2(n5003), .A3(n5004), .A4(n5005), .ZN(n4988)
         );
  NAND2_X1 U3847 ( .A1(n5006), .A2(n5007), .ZN(n5005) );
  AOI22_X1 U3848 ( .A1(n5617), .A2(n396), .B1(n5614), .B2(n6192), .ZN(n5007)
         );
  AOI22_X1 U3849 ( .A1(n5611), .A2(n6291), .B1(n5458), .B2(OUT2[11]), .ZN(
        n5006) );
  NAND2_X1 U3850 ( .A1(n5008), .A2(n5009), .ZN(n5004) );
  AOI22_X1 U3851 ( .A1(n5608), .A2(n428), .B1(n5605), .B2(n6128), .ZN(n5009)
         );
  AOI22_X1 U3852 ( .A1(n5602), .A2(n6224), .B1(n5598), .B2(n556), .ZN(n5008)
         );
  NAND2_X1 U3853 ( .A1(n5010), .A2(n5011), .ZN(n5003) );
  AOI22_X1 U3854 ( .A1(n5596), .A2(n684), .B1(n5591), .B2(n652), .ZN(n5011) );
  AOI22_X1 U3855 ( .A1(n5590), .A2(n716), .B1(n5587), .B2(n588), .ZN(n5010) );
  NAND2_X1 U3856 ( .A1(n5012), .A2(n5013), .ZN(n5002) );
  AOI22_X1 U3857 ( .A1(n5584), .A2(n492), .B1(n5581), .B2(n364), .ZN(n5013) );
  AOI22_X1 U3858 ( .A1(n5578), .A2(n524), .B1(n5573), .B2(n332), .ZN(n5012) );
  NAND2_X1 U3859 ( .A1(n5014), .A2(n5015), .ZN(n3176) );
  NOR4_X1 U3860 ( .A1(n5016), .A2(n5017), .A3(n5018), .A4(n5019), .ZN(n5015)
         );
  OAI21_X1 U3861 ( .B1(n1444), .B2(n4442), .A(n5020), .ZN(n5019) );
  NAND2_X1 U3862 ( .A1(n5664), .A2(n6473), .ZN(n5020) );
  OAI21_X1 U3863 ( .B1(n6097), .B2(n4445), .A(n5021), .ZN(n5018) );
  AOI22_X1 U3864 ( .A1(n5659), .A2(n6409), .B1(n4448), .B2(n6441), .ZN(n5021)
         );
  NAND2_X1 U3865 ( .A1(n5022), .A2(n5023), .ZN(n5017) );
  AOI22_X1 U3866 ( .A1(n5653), .A2(n2809), .B1(n4452), .B2(n6537), .ZN(n5023)
         );
  AOI22_X1 U3867 ( .A1(n5645), .A2(n6377), .B1(n4454), .B2(n6577), .ZN(n5022)
         );
  AOI22_X1 U3869 ( .A1(n5641), .A2(n6345), .B1(n4460), .B2(n6324), .ZN(n5027)
         );
  AOI22_X1 U3870 ( .A1(n5634), .A2(n6161), .B1(n4462), .B2(n6609), .ZN(n5026)
         );
  AOI22_X1 U3871 ( .A1(n5629), .A2(n2180), .B1(n4464), .B2(n6260), .ZN(n5025)
         );
  AOI22_X1 U3872 ( .A1(n4465), .A2(n619), .B1(n4466), .B2(n459), .ZN(n5024) );
  NOR4_X1 U3873 ( .A1(n5028), .A2(n5029), .A3(n5030), .A4(n5031), .ZN(n5014)
         );
  NAND2_X1 U3874 ( .A1(n5032), .A2(n5033), .ZN(n5031) );
  AOI22_X1 U3875 ( .A1(n5617), .A2(n395), .B1(n4474), .B2(n6193), .ZN(n5033)
         );
  AOI22_X1 U3876 ( .A1(n5611), .A2(n6292), .B1(n5457), .B2(OUT2[10]), .ZN(
        n5032) );
  NAND2_X1 U3877 ( .A1(n5034), .A2(n5035), .ZN(n5030) );
  AOI22_X1 U3878 ( .A1(n4478), .A2(n427), .B1(n4479), .B2(n6129), .ZN(n5035)
         );
  AOI22_X1 U3879 ( .A1(n5602), .A2(n6225), .B1(n5598), .B2(n555), .ZN(n5034)
         );
  NAND2_X1 U3880 ( .A1(n5036), .A2(n5037), .ZN(n5029) );
  AOI22_X1 U3881 ( .A1(n4484), .A2(n683), .B1(n5591), .B2(n651), .ZN(n5037) );
  AOI22_X1 U3882 ( .A1(n5590), .A2(n715), .B1(n4487), .B2(n587), .ZN(n5036) );
  NAND2_X1 U3883 ( .A1(n5038), .A2(n5039), .ZN(n5028) );
  AOI22_X1 U3884 ( .A1(n4490), .A2(n491), .B1(n4491), .B2(n363), .ZN(n5039) );
  AOI22_X1 U3885 ( .A1(n5578), .A2(n523), .B1(n5573), .B2(n331), .ZN(n5038) );
  NAND2_X1 U3886 ( .A1(n5040), .A2(n5041), .ZN(n3175) );
  NOR4_X1 U3887 ( .A1(n5042), .A2(n5043), .A3(n5044), .A4(n5045), .ZN(n5041)
         );
  OAI21_X1 U3888 ( .B1(n1445), .B2(n4442), .A(n5046), .ZN(n5045) );
  NAND2_X1 U3889 ( .A1(n5664), .A2(n6474), .ZN(n5046) );
  OAI21_X1 U3890 ( .B1(n5525), .B2(n4445), .A(n5047), .ZN(n5044) );
  AOI22_X1 U3891 ( .A1(n4447), .A2(n6410), .B1(n4448), .B2(n6442), .ZN(n5047)
         );
  NAND2_X1 U3892 ( .A1(n5048), .A2(n5049), .ZN(n5043) );
  AOI22_X1 U3893 ( .A1(n4451), .A2(n2808), .B1(n4452), .B2(n6538), .ZN(n5049)
         );
  AOI22_X1 U3894 ( .A1(n5645), .A2(n6378), .B1(n4454), .B2(n6578), .ZN(n5048)
         );
  AOI22_X1 U3896 ( .A1(n4459), .A2(n6346), .B1(n4460), .B2(n6325), .ZN(n5053)
         );
  AOI22_X1 U3897 ( .A1(n5634), .A2(n6162), .B1(n4462), .B2(n6610), .ZN(n5052)
         );
  AOI22_X1 U3898 ( .A1(n4463), .A2(n2175), .B1(n4464), .B2(n6261), .ZN(n5051)
         );
  AOI22_X1 U3899 ( .A1(n5623), .A2(n618), .B1(n4466), .B2(n458), .ZN(n5050) );
  NOR4_X1 U3900 ( .A1(n5054), .A2(n5055), .A3(n5056), .A4(n5057), .ZN(n5040)
         );
  NAND2_X1 U3901 ( .A1(n5058), .A2(n5059), .ZN(n5057) );
  AOI22_X1 U3902 ( .A1(n4473), .A2(n394), .B1(n4474), .B2(n6194), .ZN(n5059)
         );
  AOI22_X1 U3903 ( .A1(n4475), .A2(n6293), .B1(n5458), .B2(OUT2[9]), .ZN(n5058) );
  NAND2_X1 U3904 ( .A1(n5060), .A2(n5061), .ZN(n5056) );
  AOI22_X1 U3905 ( .A1(n5608), .A2(n426), .B1(n4479), .B2(n6130), .ZN(n5061)
         );
  AOI22_X1 U3906 ( .A1(n4480), .A2(n6226), .B1(n5598), .B2(n554), .ZN(n5060)
         );
  NAND2_X1 U3907 ( .A1(n5062), .A2(n5063), .ZN(n5055) );
  AOI22_X1 U3908 ( .A1(n5596), .A2(n682), .B1(n5591), .B2(n650), .ZN(n5063) );
  AOI22_X1 U3909 ( .A1(n4486), .A2(n714), .B1(n4487), .B2(n586), .ZN(n5062) );
  NAND2_X1 U3910 ( .A1(n5064), .A2(n5065), .ZN(n5054) );
  AOI22_X1 U3911 ( .A1(n5584), .A2(n490), .B1(n4491), .B2(n362), .ZN(n5065) );
  AOI22_X1 U3912 ( .A1(n4492), .A2(n522), .B1(n5573), .B2(n330), .ZN(n5064) );
  NAND2_X1 U3913 ( .A1(n5066), .A2(n5067), .ZN(n3174) );
  NOR4_X1 U3914 ( .A1(n5068), .A2(n5069), .A3(n5070), .A4(n5071), .ZN(n5067)
         );
  OAI21_X1 U3915 ( .B1(n1446), .B2(n4442), .A(n5072), .ZN(n5071) );
  NAND2_X1 U3916 ( .A1(n5664), .A2(n6475), .ZN(n5072) );
  OAI21_X1 U3917 ( .B1(n6099), .B2(n4445), .A(n5073), .ZN(n5070) );
  AOI22_X1 U3918 ( .A1(n4447), .A2(n6411), .B1(n4448), .B2(n6443), .ZN(n5073)
         );
  NAND2_X1 U3919 ( .A1(n5074), .A2(n5075), .ZN(n5069) );
  AOI22_X1 U3920 ( .A1(n4451), .A2(n2807), .B1(n4452), .B2(n6539), .ZN(n5075)
         );
  AOI22_X1 U3921 ( .A1(n5645), .A2(n6379), .B1(n4454), .B2(n6579), .ZN(n5074)
         );
  AOI22_X1 U3923 ( .A1(n4459), .A2(n6347), .B1(n4460), .B2(n6326), .ZN(n5079)
         );
  AOI22_X1 U3924 ( .A1(n5634), .A2(n6163), .B1(n4462), .B2(n6611), .ZN(n5078)
         );
  AOI22_X1 U3925 ( .A1(n4463), .A2(n2170), .B1(n4464), .B2(n6262), .ZN(n5077)
         );
  AOI22_X1 U3926 ( .A1(n4465), .A2(n617), .B1(n4466), .B2(n457), .ZN(n5076) );
  NOR4_X1 U3927 ( .A1(n5080), .A2(n5081), .A3(n5082), .A4(n5083), .ZN(n5066)
         );
  NAND2_X1 U3928 ( .A1(n5084), .A2(n5085), .ZN(n5083) );
  AOI22_X1 U3929 ( .A1(n4473), .A2(n393), .B1(n4474), .B2(n6195), .ZN(n5085)
         );
  AOI22_X1 U3930 ( .A1(n4475), .A2(n6294), .B1(n5457), .B2(OUT2[8]), .ZN(n5084) );
  NAND2_X1 U3931 ( .A1(n5086), .A2(n5087), .ZN(n5082) );
  AOI22_X1 U3932 ( .A1(n4478), .A2(n425), .B1(n4479), .B2(n6131), .ZN(n5087)
         );
  AOI22_X1 U3933 ( .A1(n4480), .A2(n6227), .B1(n5598), .B2(n553), .ZN(n5086)
         );
  NAND2_X1 U3934 ( .A1(n5088), .A2(n5089), .ZN(n5081) );
  AOI22_X1 U3935 ( .A1(n4484), .A2(n681), .B1(n5591), .B2(n649), .ZN(n5089) );
  AOI22_X1 U3936 ( .A1(n4486), .A2(n713), .B1(n4487), .B2(n585), .ZN(n5088) );
  NAND2_X1 U3937 ( .A1(n5090), .A2(n5091), .ZN(n5080) );
  AOI22_X1 U3938 ( .A1(n4490), .A2(n489), .B1(n4491), .B2(n361), .ZN(n5091) );
  AOI22_X1 U3939 ( .A1(n4492), .A2(n521), .B1(n5573), .B2(n329), .ZN(n5090) );
  NAND2_X1 U3940 ( .A1(n5092), .A2(n5093), .ZN(n3173) );
  NOR4_X1 U3941 ( .A1(n5094), .A2(n5095), .A3(n5096), .A4(n5097), .ZN(n5093)
         );
  OAI21_X1 U3942 ( .B1(n1447), .B2(n4442), .A(n5098), .ZN(n5097) );
  NAND2_X1 U3943 ( .A1(n5664), .A2(n6476), .ZN(n5098) );
  OAI21_X1 U3944 ( .B1(n6100), .B2(n4445), .A(n5099), .ZN(n5096) );
  AOI22_X1 U3945 ( .A1(n4447), .A2(n6412), .B1(n4448), .B2(n6444), .ZN(n5099)
         );
  NAND2_X1 U3946 ( .A1(n5100), .A2(n5101), .ZN(n5095) );
  AOI22_X1 U3947 ( .A1(n4451), .A2(n6548), .B1(n4452), .B2(n6540), .ZN(n5101)
         );
  AOI22_X1 U3948 ( .A1(n5645), .A2(n6380), .B1(n4454), .B2(n6580), .ZN(n5100)
         );
  AOI22_X1 U3950 ( .A1(n4459), .A2(n6348), .B1(n4460), .B2(n6327), .ZN(n5105)
         );
  AOI22_X1 U3951 ( .A1(n5634), .A2(n6164), .B1(n4462), .B2(n6612), .ZN(n5104)
         );
  AOI22_X1 U3952 ( .A1(n4463), .A2(n2165), .B1(n4464), .B2(n6263), .ZN(n5103)
         );
  AOI22_X1 U3953 ( .A1(n4465), .A2(n616), .B1(n4466), .B2(n456), .ZN(n5102) );
  NOR4_X1 U3954 ( .A1(n5106), .A2(n5107), .A3(n5108), .A4(n5109), .ZN(n5092)
         );
  NAND2_X1 U3955 ( .A1(n5110), .A2(n5111), .ZN(n5109) );
  AOI22_X1 U3956 ( .A1(n4473), .A2(n392), .B1(n4474), .B2(n6196), .ZN(n5111)
         );
  AOI22_X1 U3957 ( .A1(n4475), .A2(n6295), .B1(n5458), .B2(OUT2[7]), .ZN(n5110) );
  NAND2_X1 U3958 ( .A1(n5112), .A2(n5113), .ZN(n5108) );
  AOI22_X1 U3959 ( .A1(n4478), .A2(n424), .B1(n4479), .B2(n6132), .ZN(n5113)
         );
  AOI22_X1 U3960 ( .A1(n4480), .A2(n6228), .B1(n5598), .B2(n552), .ZN(n5112)
         );
  NAND2_X1 U3961 ( .A1(n5114), .A2(n5115), .ZN(n5107) );
  AOI22_X1 U3962 ( .A1(n4484), .A2(n680), .B1(n5591), .B2(n648), .ZN(n5115) );
  AOI22_X1 U3963 ( .A1(n4486), .A2(n712), .B1(n4487), .B2(n584), .ZN(n5114) );
  NAND2_X1 U3964 ( .A1(n5116), .A2(n5117), .ZN(n5106) );
  AOI22_X1 U3965 ( .A1(n4490), .A2(n488), .B1(n4491), .B2(n360), .ZN(n5117) );
  AOI22_X1 U3966 ( .A1(n4492), .A2(n520), .B1(n5573), .B2(n328), .ZN(n5116) );
  NAND2_X1 U3967 ( .A1(n5118), .A2(n5119), .ZN(n3172) );
  NOR4_X1 U3968 ( .A1(n5120), .A2(n5121), .A3(n5122), .A4(n5123), .ZN(n5119)
         );
  OAI21_X1 U3969 ( .B1(n1448), .B2(n4442), .A(n5124), .ZN(n5123) );
  NAND2_X1 U3970 ( .A1(n5664), .A2(n6477), .ZN(n5124) );
  OAI21_X1 U3971 ( .B1(n6101), .B2(n4445), .A(n5125), .ZN(n5122) );
  AOI22_X1 U3972 ( .A1(n4447), .A2(n6413), .B1(n4448), .B2(n6445), .ZN(n5125)
         );
  NAND2_X1 U3973 ( .A1(n5126), .A2(n5127), .ZN(n5121) );
  AOI22_X1 U3974 ( .A1(n4451), .A2(n6549), .B1(n4452), .B2(n6541), .ZN(n5127)
         );
  AOI22_X1 U3975 ( .A1(n5645), .A2(n6381), .B1(n4454), .B2(n6581), .ZN(n5126)
         );
  AOI22_X1 U3977 ( .A1(n4459), .A2(n6349), .B1(n4460), .B2(n6328), .ZN(n5131)
         );
  AOI22_X1 U3978 ( .A1(n5634), .A2(n6165), .B1(n4462), .B2(n6613), .ZN(n5130)
         );
  AOI22_X1 U3979 ( .A1(n4463), .A2(n2160), .B1(n4464), .B2(n6264), .ZN(n5129)
         );
  AOI22_X1 U3980 ( .A1(n4465), .A2(n615), .B1(n4466), .B2(n455), .ZN(n5128) );
  NOR4_X1 U3981 ( .A1(n5132), .A2(n5133), .A3(n5134), .A4(n5135), .ZN(n5118)
         );
  NAND2_X1 U3982 ( .A1(n5136), .A2(n5137), .ZN(n5135) );
  AOI22_X1 U3983 ( .A1(n4473), .A2(n391), .B1(n4474), .B2(n6197), .ZN(n5137)
         );
  AOI22_X1 U3984 ( .A1(n4475), .A2(n6296), .B1(n5457), .B2(OUT2[6]), .ZN(n5136) );
  NAND2_X1 U3985 ( .A1(n5138), .A2(n5139), .ZN(n5134) );
  AOI22_X1 U3986 ( .A1(n4478), .A2(n423), .B1(n4479), .B2(n6133), .ZN(n5139)
         );
  AOI22_X1 U3987 ( .A1(n4480), .A2(n6229), .B1(n5598), .B2(n551), .ZN(n5138)
         );
  NAND2_X1 U3988 ( .A1(n5140), .A2(n5141), .ZN(n5133) );
  AOI22_X1 U3989 ( .A1(n4484), .A2(n679), .B1(n5591), .B2(n647), .ZN(n5141) );
  AOI22_X1 U3990 ( .A1(n4486), .A2(n711), .B1(n4487), .B2(n583), .ZN(n5140) );
  NAND2_X1 U3991 ( .A1(n5142), .A2(n5143), .ZN(n5132) );
  AOI22_X1 U3992 ( .A1(n4490), .A2(n487), .B1(n4491), .B2(n359), .ZN(n5143) );
  AOI22_X1 U3993 ( .A1(n4492), .A2(n519), .B1(n5573), .B2(n327), .ZN(n5142) );
  NAND2_X1 U3994 ( .A1(n5144), .A2(n5145), .ZN(n3171) );
  NOR4_X1 U3995 ( .A1(n5146), .A2(n5147), .A3(n5148), .A4(n5149), .ZN(n5145)
         );
  OAI21_X1 U3996 ( .B1(n1449), .B2(n4442), .A(n5150), .ZN(n5149) );
  NAND2_X1 U3997 ( .A1(n5664), .A2(n6478), .ZN(n5150) );
  OAI21_X1 U3998 ( .B1(n6102), .B2(n4445), .A(n5151), .ZN(n5148) );
  AOI22_X1 U3999 ( .A1(n4447), .A2(n6414), .B1(n4448), .B2(n6446), .ZN(n5151)
         );
  NAND2_X1 U4000 ( .A1(n5152), .A2(n5153), .ZN(n5147) );
  AOI22_X1 U4001 ( .A1(n4451), .A2(n6550), .B1(n4452), .B2(n6542), .ZN(n5153)
         );
  AOI22_X1 U4002 ( .A1(n5645), .A2(n6382), .B1(n4454), .B2(n6582), .ZN(n5152)
         );
  AOI22_X1 U4004 ( .A1(n4459), .A2(n6350), .B1(n4460), .B2(n6329), .ZN(n5157)
         );
  AOI22_X1 U4005 ( .A1(n5634), .A2(n6166), .B1(n4462), .B2(n6614), .ZN(n5156)
         );
  AOI22_X1 U4006 ( .A1(n4463), .A2(n2155), .B1(n4464), .B2(n6265), .ZN(n5155)
         );
  AOI22_X1 U4007 ( .A1(n4465), .A2(n614), .B1(n4466), .B2(n454), .ZN(n5154) );
  NOR4_X1 U4008 ( .A1(n5158), .A2(n5159), .A3(n5160), .A4(n5161), .ZN(n5144)
         );
  NAND2_X1 U4009 ( .A1(n5162), .A2(n5163), .ZN(n5161) );
  AOI22_X1 U4010 ( .A1(n4473), .A2(n390), .B1(n4474), .B2(n6198), .ZN(n5163)
         );
  AOI22_X1 U4011 ( .A1(n4475), .A2(n6297), .B1(n5458), .B2(OUT2[5]), .ZN(n5162) );
  NAND2_X1 U4012 ( .A1(n5164), .A2(n5165), .ZN(n5160) );
  AOI22_X1 U4013 ( .A1(n4478), .A2(n422), .B1(n4479), .B2(n6134), .ZN(n5165)
         );
  AOI22_X1 U4014 ( .A1(n4480), .A2(n6230), .B1(n5598), .B2(n550), .ZN(n5164)
         );
  NAND2_X1 U4015 ( .A1(n5166), .A2(n5167), .ZN(n5159) );
  AOI22_X1 U4016 ( .A1(n4484), .A2(n678), .B1(n5591), .B2(n646), .ZN(n5167) );
  AOI22_X1 U4017 ( .A1(n4486), .A2(n710), .B1(n4487), .B2(n582), .ZN(n5166) );
  NAND2_X1 U4018 ( .A1(n5168), .A2(n5169), .ZN(n5158) );
  AOI22_X1 U4019 ( .A1(n4490), .A2(n486), .B1(n4491), .B2(n358), .ZN(n5169) );
  AOI22_X1 U4020 ( .A1(n4492), .A2(n518), .B1(n5573), .B2(n326), .ZN(n5168) );
  NAND2_X1 U4021 ( .A1(n5170), .A2(n5171), .ZN(n3170) );
  NOR4_X1 U4022 ( .A1(n5172), .A2(n5173), .A3(n5174), .A4(n5175), .ZN(n5171)
         );
  OAI21_X1 U4023 ( .B1(n1450), .B2(n4442), .A(n5176), .ZN(n5175) );
  NAND2_X1 U4024 ( .A1(n5664), .A2(n6479), .ZN(n5176) );
  OAI21_X1 U4025 ( .B1(n6103), .B2(n4445), .A(n5177), .ZN(n5174) );
  AOI22_X1 U4026 ( .A1(n4447), .A2(n6415), .B1(n4448), .B2(n6447), .ZN(n5177)
         );
  NAND2_X1 U4027 ( .A1(n5178), .A2(n5179), .ZN(n5173) );
  AOI22_X1 U4028 ( .A1(n4451), .A2(n6551), .B1(n4452), .B2(n6543), .ZN(n5179)
         );
  AOI22_X1 U4029 ( .A1(n5645), .A2(n6383), .B1(n4454), .B2(n6583), .ZN(n5178)
         );
  AOI22_X1 U4031 ( .A1(n4459), .A2(n6351), .B1(n4460), .B2(n6330), .ZN(n5183)
         );
  AOI22_X1 U4032 ( .A1(n5634), .A2(n6167), .B1(n4462), .B2(n6615), .ZN(n5182)
         );
  AOI22_X1 U4033 ( .A1(n4463), .A2(n2150), .B1(n4464), .B2(n6266), .ZN(n5181)
         );
  AOI22_X1 U4034 ( .A1(n4465), .A2(n613), .B1(n4466), .B2(n453), .ZN(n5180) );
  NOR4_X1 U4035 ( .A1(n5184), .A2(n5185), .A3(n5186), .A4(n5187), .ZN(n5170)
         );
  NAND2_X1 U4036 ( .A1(n5188), .A2(n5189), .ZN(n5187) );
  AOI22_X1 U4037 ( .A1(n4473), .A2(n389), .B1(n4474), .B2(n6199), .ZN(n5189)
         );
  AOI22_X1 U4038 ( .A1(n4475), .A2(n6298), .B1(n5458), .B2(OUT2[4]), .ZN(n5188) );
  NAND2_X1 U4039 ( .A1(n5190), .A2(n5191), .ZN(n5186) );
  AOI22_X1 U4040 ( .A1(n4478), .A2(n421), .B1(n4479), .B2(n6135), .ZN(n5191)
         );
  AOI22_X1 U4041 ( .A1(n4480), .A2(n6231), .B1(n5598), .B2(n549), .ZN(n5190)
         );
  NAND2_X1 U4042 ( .A1(n5192), .A2(n5193), .ZN(n5185) );
  AOI22_X1 U4043 ( .A1(n4484), .A2(n677), .B1(n5591), .B2(n645), .ZN(n5193) );
  AOI22_X1 U4044 ( .A1(n4486), .A2(n709), .B1(n4487), .B2(n581), .ZN(n5192) );
  NAND2_X1 U4045 ( .A1(n5194), .A2(n5195), .ZN(n5184) );
  AOI22_X1 U4046 ( .A1(n4490), .A2(n485), .B1(n4491), .B2(n357), .ZN(n5195) );
  AOI22_X1 U4047 ( .A1(n4492), .A2(n517), .B1(n5573), .B2(n325), .ZN(n5194) );
  NAND2_X1 U4048 ( .A1(n5196), .A2(n5197), .ZN(n3169) );
  NOR4_X1 U4049 ( .A1(n5198), .A2(n5199), .A3(n5200), .A4(n5201), .ZN(n5197)
         );
  OAI21_X1 U4050 ( .B1(n1451), .B2(n4442), .A(n5202), .ZN(n5201) );
  NAND2_X1 U4051 ( .A1(n5664), .A2(n6480), .ZN(n5202) );
  OAI21_X1 U4052 ( .B1(n6104), .B2(n4445), .A(n5203), .ZN(n5200) );
  AOI22_X1 U4053 ( .A1(n4447), .A2(n6416), .B1(n4448), .B2(n6448), .ZN(n5203)
         );
  NAND2_X1 U4054 ( .A1(n5204), .A2(n5205), .ZN(n5199) );
  AOI22_X1 U4055 ( .A1(n4451), .A2(n6552), .B1(n4452), .B2(n6544), .ZN(n5205)
         );
  AOI22_X1 U4056 ( .A1(n5645), .A2(n6384), .B1(n4454), .B2(n6584), .ZN(n5204)
         );
  AOI22_X1 U4058 ( .A1(n4459), .A2(n6352), .B1(n4460), .B2(n6331), .ZN(n5209)
         );
  AOI22_X1 U4059 ( .A1(n5634), .A2(n6168), .B1(n4462), .B2(n6616), .ZN(n5208)
         );
  AOI22_X1 U4060 ( .A1(n4463), .A2(n2145), .B1(n4464), .B2(n6267), .ZN(n5207)
         );
  AOI22_X1 U4061 ( .A1(n4465), .A2(n612), .B1(n4466), .B2(n452), .ZN(n5206) );
  NOR4_X1 U4062 ( .A1(n5210), .A2(n5211), .A3(n5212), .A4(n5213), .ZN(n5196)
         );
  NAND2_X1 U4063 ( .A1(n5214), .A2(n5215), .ZN(n5213) );
  AOI22_X1 U4064 ( .A1(n5617), .A2(n388), .B1(n5614), .B2(n6200), .ZN(n5215)
         );
  AOI22_X1 U4065 ( .A1(n5611), .A2(n6299), .B1(n5458), .B2(OUT2[3]), .ZN(n5214) );
  NAND2_X1 U4066 ( .A1(n5216), .A2(n5217), .ZN(n5212) );
  AOI22_X1 U4067 ( .A1(n4478), .A2(n420), .B1(n4479), .B2(n6136), .ZN(n5217)
         );
  AOI22_X1 U4068 ( .A1(n4480), .A2(n6232), .B1(n5598), .B2(n548), .ZN(n5216)
         );
  NAND2_X1 U4069 ( .A1(n5218), .A2(n5219), .ZN(n5211) );
  AOI22_X1 U4070 ( .A1(n4484), .A2(n676), .B1(n5591), .B2(n644), .ZN(n5219) );
  AOI22_X1 U4071 ( .A1(n4486), .A2(n708), .B1(n4487), .B2(n580), .ZN(n5218) );
  NAND2_X1 U4072 ( .A1(n5220), .A2(n5221), .ZN(n5210) );
  AOI22_X1 U4073 ( .A1(n4490), .A2(n484), .B1(n4491), .B2(n356), .ZN(n5221) );
  AOI22_X1 U4074 ( .A1(n4492), .A2(n516), .B1(n5573), .B2(n324), .ZN(n5220) );
  NAND2_X1 U4075 ( .A1(n5222), .A2(n5223), .ZN(n3168) );
  NOR4_X1 U4076 ( .A1(n5224), .A2(n5225), .A3(n5226), .A4(n5227), .ZN(n5223)
         );
  OAI21_X1 U4077 ( .B1(n1452), .B2(n4442), .A(n5228), .ZN(n5227) );
  NAND2_X1 U4078 ( .A1(n5664), .A2(n6481), .ZN(n5228) );
  OAI21_X1 U4079 ( .B1(n6105), .B2(n4445), .A(n5229), .ZN(n5226) );
  AOI22_X1 U4080 ( .A1(n4447), .A2(n6417), .B1(n4448), .B2(n6449), .ZN(n5229)
         );
  NAND2_X1 U4081 ( .A1(n5230), .A2(n5231), .ZN(n5225) );
  AOI22_X1 U4082 ( .A1(n4451), .A2(n6553), .B1(n4452), .B2(n6545), .ZN(n5231)
         );
  AOI22_X1 U4083 ( .A1(n5645), .A2(n6385), .B1(n4454), .B2(n6585), .ZN(n5230)
         );
  AOI22_X1 U4085 ( .A1(n4459), .A2(n6353), .B1(n4460), .B2(n6332), .ZN(n5235)
         );
  AOI22_X1 U4086 ( .A1(n5634), .A2(n6169), .B1(n4462), .B2(n6617), .ZN(n5234)
         );
  AOI22_X1 U4087 ( .A1(n4463), .A2(n2140), .B1(n4464), .B2(n6268), .ZN(n5233)
         );
  AOI22_X1 U4088 ( .A1(n4465), .A2(n611), .B1(n4466), .B2(n451), .ZN(n5232) );
  NOR4_X1 U4089 ( .A1(n5236), .A2(n5237), .A3(n5238), .A4(n5239), .ZN(n5222)
         );
  NAND2_X1 U4090 ( .A1(n5240), .A2(n5241), .ZN(n5239) );
  AOI22_X1 U4091 ( .A1(n4473), .A2(n387), .B1(n4474), .B2(n6201), .ZN(n5241)
         );
  AOI22_X1 U4092 ( .A1(n4475), .A2(n6300), .B1(n5457), .B2(OUT2[2]), .ZN(n5240) );
  NAND2_X1 U4093 ( .A1(n5242), .A2(n5243), .ZN(n5238) );
  AOI22_X1 U4094 ( .A1(n4478), .A2(n419), .B1(n4479), .B2(n6137), .ZN(n5243)
         );
  AOI22_X1 U4095 ( .A1(n4480), .A2(n6233), .B1(n5598), .B2(n547), .ZN(n5242)
         );
  NAND2_X1 U4096 ( .A1(n5244), .A2(n5245), .ZN(n5237) );
  AOI22_X1 U4097 ( .A1(n4484), .A2(n675), .B1(n5591), .B2(n643), .ZN(n5245) );
  AOI22_X1 U4098 ( .A1(n4486), .A2(n707), .B1(n4487), .B2(n579), .ZN(n5244) );
  NAND2_X1 U4099 ( .A1(n5246), .A2(n5247), .ZN(n5236) );
  AOI22_X1 U4100 ( .A1(n4490), .A2(n483), .B1(n4491), .B2(n355), .ZN(n5247) );
  AOI22_X1 U4101 ( .A1(n4492), .A2(n515), .B1(n5573), .B2(n323), .ZN(n5246) );
  NAND2_X1 U4102 ( .A1(n5248), .A2(n5249), .ZN(n3167) );
  NOR4_X1 U4103 ( .A1(n5250), .A2(n5251), .A3(n5252), .A4(n5253), .ZN(n5249)
         );
  OAI21_X1 U4104 ( .B1(n1453), .B2(n4442), .A(n5254), .ZN(n5253) );
  NAND2_X1 U4105 ( .A1(n5664), .A2(n6482), .ZN(n5254) );
  OAI21_X1 U4106 ( .B1(n6106), .B2(n4445), .A(n5255), .ZN(n5252) );
  AOI22_X1 U4107 ( .A1(n4447), .A2(n6418), .B1(n4448), .B2(n6450), .ZN(n5255)
         );
  NAND2_X1 U4108 ( .A1(n5256), .A2(n5257), .ZN(n5251) );
  AOI22_X1 U4109 ( .A1(n4451), .A2(n6554), .B1(n4452), .B2(n6546), .ZN(n5257)
         );
  AOI22_X1 U4110 ( .A1(n5645), .A2(n6386), .B1(n4454), .B2(n6586), .ZN(n5256)
         );
  AOI22_X1 U4112 ( .A1(n4459), .A2(n6354), .B1(n4460), .B2(n6333), .ZN(n5261)
         );
  AOI22_X1 U4113 ( .A1(n4461), .A2(n6170), .B1(n4462), .B2(n6618), .ZN(n5260)
         );
  AOI22_X1 U4114 ( .A1(n4463), .A2(n2135), .B1(n4464), .B2(n6269), .ZN(n5259)
         );
  AOI22_X1 U4115 ( .A1(n4465), .A2(n610), .B1(n4466), .B2(n450), .ZN(n5258) );
  NOR4_X1 U4116 ( .A1(n5262), .A2(n5263), .A3(n5264), .A4(n5265), .ZN(n5248)
         );
  NAND2_X1 U4117 ( .A1(n5266), .A2(n5267), .ZN(n5265) );
  AOI22_X1 U4118 ( .A1(n4473), .A2(n386), .B1(n4474), .B2(n6202), .ZN(n5267)
         );
  AOI22_X1 U4119 ( .A1(n4475), .A2(n6301), .B1(n5457), .B2(OUT2[1]), .ZN(n5266) );
  NAND2_X1 U4120 ( .A1(n5268), .A2(n5269), .ZN(n5264) );
  AOI22_X1 U4121 ( .A1(n4478), .A2(n418), .B1(n4479), .B2(n6138), .ZN(n5269)
         );
  AOI22_X1 U4122 ( .A1(n4480), .A2(n6234), .B1(n5598), .B2(n546), .ZN(n5268)
         );
  NAND2_X1 U4123 ( .A1(n5270), .A2(n5271), .ZN(n5263) );
  AOI22_X1 U4124 ( .A1(n4484), .A2(n674), .B1(n5591), .B2(n642), .ZN(n5271) );
  AOI22_X1 U4125 ( .A1(n4486), .A2(n706), .B1(n4487), .B2(n578), .ZN(n5270) );
  NAND2_X1 U4126 ( .A1(n5272), .A2(n5273), .ZN(n5262) );
  AOI22_X1 U4127 ( .A1(n4490), .A2(n482), .B1(n4491), .B2(n354), .ZN(n5273) );
  AOI22_X1 U4128 ( .A1(n4492), .A2(n514), .B1(n5573), .B2(n322), .ZN(n5272) );
  NAND2_X1 U4129 ( .A1(n5274), .A2(n5275), .ZN(n3166) );
  NOR4_X1 U4130 ( .A1(n5276), .A2(n5277), .A3(n5278), .A4(n5279), .ZN(n5275)
         );
  OAI21_X1 U4131 ( .B1(n1454), .B2(n5668), .A(n5280), .ZN(n5279) );
  NAND2_X1 U4132 ( .A1(n5664), .A2(n6483), .ZN(n5280) );
  NOR2_X1 U4133 ( .A1(n5281), .A2(n5282), .ZN(n4444) );
  OR2_X1 U4134 ( .A1(n5281), .A2(n5283), .ZN(n4442) );
  OAI21_X1 U4135 ( .B1(n6107), .B2(n5662), .A(n5284), .ZN(n5278) );
  AOI22_X1 U4136 ( .A1(n5659), .A2(n6419), .B1(n5656), .B2(n6451), .ZN(n5284)
         );
  NOR2_X1 U4137 ( .A1(n5283), .A2(n5285), .ZN(n4448) );
  NOR2_X1 U4138 ( .A1(n5285), .A2(n5282), .ZN(n4447) );
  NAND2_X1 U4139 ( .A1(n5286), .A2(n5287), .ZN(n4445) );
  NOR4_X1 U4140 ( .A1(n6620), .A2(n5288), .A3(n5289), .A4(n5290), .ZN(n5287)
         );
  NOR3_X1 U4141 ( .A1(n5291), .A2(n5292), .A3(n5293), .ZN(n5286) );
  NAND2_X1 U4142 ( .A1(n5294), .A2(n5295), .ZN(n5277) );
  AOI22_X1 U4143 ( .A1(n5653), .A2(n6555), .B1(n5650), .B2(n6547), .ZN(n5295)
         );
  NOR2_X1 U4144 ( .A1(n5296), .A2(n5297), .ZN(n4452) );
  NOR2_X1 U4145 ( .A1(n5297), .A2(n5298), .ZN(n4451) );
  AOI22_X1 U4146 ( .A1(n5645), .A2(n6387), .B1(n5644), .B2(n6587), .ZN(n5294)
         );
  NOR2_X1 U4147 ( .A1(n5299), .A2(n5296), .ZN(n4454) );
  NOR2_X1 U4148 ( .A1(n5297), .A2(n5283), .ZN(n4453) );
  AOI22_X1 U4150 ( .A1(n5641), .A2(n6355), .B1(n5638), .B2(n6334), .ZN(n5303)
         );
  NOR2_X1 U4151 ( .A1(n5304), .A2(n5281), .ZN(n4460) );
  NOR2_X1 U4152 ( .A1(n5305), .A2(n5281), .ZN(n4459) );
  AOI22_X1 U4153 ( .A1(n5634), .A2(n6171), .B1(n5632), .B2(n6619), .ZN(n5302)
         );
  NOR2_X1 U4154 ( .A1(n5299), .A2(n5298), .ZN(n4462) );
  NOR2_X1 U4155 ( .A1(n5299), .A2(n5306), .ZN(n4461) );
  AOI22_X1 U4156 ( .A1(n5629), .A2(n2130), .B1(n5626), .B2(n6270), .ZN(n5301)
         );
  NOR2_X1 U4157 ( .A1(n5305), .A2(n5285), .ZN(n4464) );
  NOR2_X1 U4158 ( .A1(n5304), .A2(n5285), .ZN(n4463) );
  AOI22_X1 U4159 ( .A1(n5623), .A2(n609), .B1(n5620), .B2(n449), .ZN(n5300) );
  NOR2_X1 U4160 ( .A1(n5307), .A2(n5281), .ZN(n4466) );
  NOR2_X1 U4161 ( .A1(n5307), .A2(n5297), .ZN(n4465) );
  NOR4_X1 U4162 ( .A1(n5308), .A2(n5309), .A3(n5310), .A4(n5311), .ZN(n5274)
         );
  NAND2_X1 U4163 ( .A1(n5312), .A2(n5313), .ZN(n5311) );
  AOI22_X1 U4164 ( .A1(n4473), .A2(n385), .B1(n4474), .B2(n6203), .ZN(n5313)
         );
  NOR2_X1 U4165 ( .A1(n5307), .A2(n5299), .ZN(n4474) );
  NOR2_X1 U4166 ( .A1(n5304), .A2(n5299), .ZN(n4473) );
  AOI22_X1 U4167 ( .A1(n4475), .A2(n6302), .B1(n5457), .B2(OUT2[0]), .ZN(n5312) );
  NOR2_X1 U4168 ( .A1(n5305), .A2(n5299), .ZN(n4475) );
  NAND2_X1 U4169 ( .A1(n5314), .A2(n5315), .ZN(n5310) );
  AOI22_X1 U4170 ( .A1(n5608), .A2(n417), .B1(n5605), .B2(n6139), .ZN(n5315)
         );
  NOR2_X1 U4171 ( .A1(n5285), .A2(n5306), .ZN(n4479) );
  NOR2_X1 U4172 ( .A1(n5305), .A2(n5297), .ZN(n4478) );
  NAND2_X1 U4173 ( .A1(n5316), .A2(ADD_RD2[3]), .ZN(n5305) );
  NOR2_X1 U4174 ( .A1(ADD_RD2[4]), .A2(n6075), .ZN(n5316) );
  AOI22_X1 U4175 ( .A1(n5602), .A2(n6235), .B1(n5598), .B2(n545), .ZN(n5314)
         );
  NOR2_X1 U4176 ( .A1(n5304), .A2(n5297), .ZN(n4481) );
  NAND2_X1 U4177 ( .A1(n5317), .A2(ADD_RD2[3]), .ZN(n5304) );
  NOR2_X1 U4178 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[0]), .ZN(n5317) );
  NOR2_X1 U4179 ( .A1(n5281), .A2(n5306), .ZN(n4480) );
  NAND2_X1 U4180 ( .A1(n5318), .A2(n5319), .ZN(n5309) );
  AOI22_X1 U4181 ( .A1(n5596), .A2(n673), .B1(n5591), .B2(n641), .ZN(n5319) );
  NOR2_X1 U4182 ( .A1(n5298), .A2(n5285), .ZN(n4485) );
  NOR2_X1 U4183 ( .A1(n5297), .A2(n5282), .ZN(n4484) );
  NAND2_X1 U4184 ( .A1(n5320), .A2(n5321), .ZN(n5297) );
  NOR2_X1 U4185 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n5320) );
  AOI22_X1 U4186 ( .A1(n5590), .A2(n705), .B1(n5587), .B2(n577), .ZN(n5318) );
  NOR2_X1 U4187 ( .A1(n5307), .A2(n5285), .ZN(n4487) );
  OR2_X1 U4188 ( .A1(n5322), .A2(n6075), .ZN(n5307) );
  OR2_X1 U4189 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n5322) );
  NOR2_X1 U4190 ( .A1(n5299), .A2(n5282), .ZN(n4486) );
  OR2_X1 U4191 ( .A1(n5323), .A2(n6072), .ZN(n5282) );
  OR2_X1 U4192 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[0]), .ZN(n5323) );
  NAND2_X1 U4193 ( .A1(n5324), .A2(n5325), .ZN(n5308) );
  AOI22_X1 U4194 ( .A1(n5584), .A2(n481), .B1(n5581), .B2(n353), .ZN(n5325) );
  NOR2_X1 U4195 ( .A1(n5296), .A2(n5281), .ZN(n4491) );
  NOR2_X1 U4196 ( .A1(n5296), .A2(n5285), .ZN(n4490) );
  NAND2_X1 U4197 ( .A1(n5326), .A2(n5321), .ZN(n5285) );
  NOR2_X1 U4198 ( .A1(ADD_RD2[2]), .A2(n6074), .ZN(n5326) );
  NAND2_X1 U4199 ( .A1(n5327), .A2(ADD_RD2[3]), .ZN(n5296) );
  NOR2_X1 U4200 ( .A1(ADD_RD2[0]), .A2(n6072), .ZN(n5327) );
  AOI22_X1 U4201 ( .A1(n5578), .A2(n513), .B1(n5573), .B2(n321), .ZN(n5324) );
  NOR2_X1 U4202 ( .A1(n5298), .A2(n5281), .ZN(n4493) );
  NAND2_X1 U4203 ( .A1(n5328), .A2(n5321), .ZN(n5281) );
  NOR2_X1 U4204 ( .A1(n6073), .A2(n6074), .ZN(n5328) );
  NAND2_X1 U4205 ( .A1(n5329), .A2(ADD_RD2[3]), .ZN(n5298) );
  NOR2_X1 U4206 ( .A1(n6072), .A2(n6075), .ZN(n5329) );
  NOR2_X1 U4207 ( .A1(n5299), .A2(n5283), .ZN(n4492) );
  OR2_X1 U4208 ( .A1(n5330), .A2(n6075), .ZN(n5283) );
  OR2_X1 U4209 ( .A1(ADD_RD2[3]), .A2(n6072), .ZN(n5330) );
  NAND2_X1 U4210 ( .A1(n5331), .A2(n5321), .ZN(n5299) );
  NOR2_X1 U4211 ( .A1(n5291), .A2(n5332), .ZN(n5321) );
  XOR2_X1 U4214 ( .A(ADD_WR[3]), .B(ADD_RD2[3]), .Z(n5288) );
  XOR2_X1 U4215 ( .A(ADD_RD2[1]), .B(ADD_WR[1]), .Z(n5289) );
  XOR2_X1 U4217 ( .A(ADD_WR[4]), .B(ADD_RD2[4]), .Z(n5292) );
  XOR2_X1 U4218 ( .A(ADD_RD2[0]), .B(ADD_WR[0]), .Z(n5290) );
  XOR2_X1 U4219 ( .A(ADD_RD2[2]), .B(ADD_WR[2]), .Z(n5293) );
  NAND2_X1 U4220 ( .A1(n5335), .A2(RD2), .ZN(n5291) );
  NOR2_X1 U4221 ( .A1(n5336), .A2(n5939), .ZN(n5335) );
  NOR3_X1 U4222 ( .A1(n5306), .A2(ADD_RD2[2]), .A3(ADD_RD2[1]), .ZN(n5336) );
  NAND2_X1 U4223 ( .A1(n5337), .A2(n6075), .ZN(n5306) );
  NOR2_X1 U4224 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n5337) );
  NOR2_X1 U4225 ( .A1(ADD_RD2[1]), .A2(n6073), .ZN(n5331) );
  OAI21_X1 U4226 ( .B1(n6093), .B2(n1828), .A(n5338), .ZN(n3165) );
  NAND2_X1 U4227 ( .A1(n1828), .A2(n6437), .ZN(n5338) );
  OAI21_X1 U4228 ( .B1(n6094), .B2(n1828), .A(n5339), .ZN(n3164) );
  NAND2_X1 U4229 ( .A1(n5868), .A2(n6438), .ZN(n5339) );
  OAI21_X1 U4230 ( .B1(n6095), .B2(n1828), .A(n5340), .ZN(n3163) );
  NAND2_X1 U4231 ( .A1(n5868), .A2(n6439), .ZN(n5340) );
  OAI21_X1 U4232 ( .B1(n6096), .B2(n1828), .A(n5341), .ZN(n3162) );
  NAND2_X1 U4233 ( .A1(n5868), .A2(n6440), .ZN(n5341) );
  OAI21_X1 U4234 ( .B1(n6097), .B2(n1828), .A(n5342), .ZN(n3161) );
  NAND2_X1 U4235 ( .A1(n5868), .A2(n6441), .ZN(n5342) );
  OAI21_X1 U4236 ( .B1(n5525), .B2(n5872), .A(n5343), .ZN(n3160) );
  NAND2_X1 U4237 ( .A1(n5868), .A2(n6442), .ZN(n5343) );
  OAI21_X1 U4238 ( .B1(n6099), .B2(n5872), .A(n5344), .ZN(n3159) );
  NAND2_X1 U4239 ( .A1(n5868), .A2(n6443), .ZN(n5344) );
  OAI21_X1 U4240 ( .B1(n6100), .B2(n5872), .A(n5345), .ZN(n3158) );
  NAND2_X1 U4241 ( .A1(n5868), .A2(n6444), .ZN(n5345) );
  OAI21_X1 U4242 ( .B1(n6101), .B2(n5872), .A(n5346), .ZN(n3157) );
  NAND2_X1 U4243 ( .A1(n1828), .A2(n6445), .ZN(n5346) );
  OAI21_X1 U4244 ( .B1(n6102), .B2(n5872), .A(n5347), .ZN(n3156) );
  NAND2_X1 U4245 ( .A1(n1828), .A2(n6446), .ZN(n5347) );
  OAI21_X1 U4246 ( .B1(n6103), .B2(n5872), .A(n5348), .ZN(n3155) );
  NAND2_X1 U4247 ( .A1(n1828), .A2(n6447), .ZN(n5348) );
  OAI21_X1 U4248 ( .B1(n6104), .B2(n5872), .A(n5349), .ZN(n3154) );
  NAND2_X1 U4249 ( .A1(n1828), .A2(n6448), .ZN(n5349) );
  OAI21_X1 U4250 ( .B1(n6105), .B2(n5872), .A(n5350), .ZN(n3153) );
  NAND2_X1 U4251 ( .A1(n5868), .A2(n6449), .ZN(n5350) );
  OAI21_X1 U4252 ( .B1(n6106), .B2(n5872), .A(n5351), .ZN(n3152) );
  NAND2_X1 U4253 ( .A1(n1828), .A2(n6450), .ZN(n5351) );
  OAI21_X1 U4254 ( .B1(n6107), .B2(n1828), .A(n5352), .ZN(n3151) );
  NAND2_X1 U4255 ( .A1(n5872), .A2(n6451), .ZN(n5352) );
  NAND2_X1 U4256 ( .A1(n1692), .A2(n1590), .ZN(n1828) );
  NOR2_X1 U4258 ( .A1(ADD_WR[2]), .A2(n6067), .ZN(n5353) );
  NOR2_X1 U4259 ( .A1(n5354), .A2(n6064), .ZN(n1692) );
  OR2_X1 U4260 ( .A1(ADD_WR[3]), .A2(n2273), .ZN(n5354) );
  OAI21_X1 U4261 ( .B1(n6076), .B2(n5570), .A(n5356), .ZN(n3150) );
  NAND2_X1 U4262 ( .A1(n5355), .A2(n6588), .ZN(n5356) );
  OAI21_X1 U4263 ( .B1(n6077), .B2(n5570), .A(n5357), .ZN(n3149) );
  NAND2_X1 U4264 ( .A1(n5355), .A2(n6589), .ZN(n5357) );
  OAI21_X1 U4265 ( .B1(n6078), .B2(n5570), .A(n5358), .ZN(n3148) );
  NAND2_X1 U4266 ( .A1(n5355), .A2(n6590), .ZN(n5358) );
  OAI21_X1 U4267 ( .B1(n6079), .B2(n5570), .A(n5359), .ZN(n3147) );
  NAND2_X1 U4268 ( .A1(n5355), .A2(n6591), .ZN(n5359) );
  OAI21_X1 U4269 ( .B1(n6080), .B2(n5570), .A(n5360), .ZN(n3146) );
  NAND2_X1 U4270 ( .A1(n5355), .A2(n6592), .ZN(n5360) );
  OAI21_X1 U4271 ( .B1(n6081), .B2(n5570), .A(n5361), .ZN(n3145) );
  NAND2_X1 U4272 ( .A1(n5572), .A2(n6593), .ZN(n5361) );
  OAI21_X1 U4273 ( .B1(n5477), .B2(n5570), .A(n5362), .ZN(n3144) );
  NAND2_X1 U4274 ( .A1(n5572), .A2(n6594), .ZN(n5362) );
  OAI21_X1 U4275 ( .B1(n6083), .B2(n5570), .A(n5363), .ZN(n3143) );
  NAND2_X1 U4276 ( .A1(n5570), .A2(n6595), .ZN(n5363) );
  OAI21_X1 U4277 ( .B1(n6084), .B2(n5570), .A(n5364), .ZN(n3142) );
  NAND2_X1 U4278 ( .A1(n5572), .A2(n6596), .ZN(n5364) );
  OAI21_X1 U4279 ( .B1(n6085), .B2(n5570), .A(n5365), .ZN(n3141) );
  NAND2_X1 U4280 ( .A1(n5572), .A2(n6597), .ZN(n5365) );
  OAI21_X1 U4281 ( .B1(n6086), .B2(n5570), .A(n5366), .ZN(n3140) );
  NAND2_X1 U4282 ( .A1(n5570), .A2(n6598), .ZN(n5366) );
  OAI21_X1 U4283 ( .B1(n6087), .B2(n5570), .A(n5367), .ZN(n3139) );
  NAND2_X1 U4284 ( .A1(n5355), .A2(n6599), .ZN(n5367) );
  OAI21_X1 U4285 ( .B1(n6088), .B2(n5572), .A(n5368), .ZN(n3138) );
  NAND2_X1 U4286 ( .A1(n5355), .A2(n6600), .ZN(n5368) );
  OAI21_X1 U4287 ( .B1(n6089), .B2(n5570), .A(n5369), .ZN(n3137) );
  NAND2_X1 U4288 ( .A1(n5355), .A2(n6601), .ZN(n5369) );
  OAI21_X1 U4289 ( .B1(n6090), .B2(n5570), .A(n5370), .ZN(n3136) );
  NAND2_X1 U4290 ( .A1(n5355), .A2(n6602), .ZN(n5370) );
  OAI21_X1 U4291 ( .B1(n6091), .B2(n5572), .A(n5371), .ZN(n3135) );
  NAND2_X1 U4292 ( .A1(n5355), .A2(n6603), .ZN(n5371) );
  OAI21_X1 U4293 ( .B1(n5507), .B2(n5570), .A(n5372), .ZN(n3134) );
  NAND2_X1 U4294 ( .A1(n5355), .A2(n6604), .ZN(n5372) );
  OAI21_X1 U4295 ( .B1(n6093), .B2(n5572), .A(n5373), .ZN(n3133) );
  NAND2_X1 U4296 ( .A1(n5355), .A2(n6605), .ZN(n5373) );
  OAI21_X1 U4297 ( .B1(n6094), .B2(n5570), .A(n5374), .ZN(n3132) );
  NAND2_X1 U4298 ( .A1(n5355), .A2(n6606), .ZN(n5374) );
  OAI21_X1 U4299 ( .B1(n6095), .B2(n5572), .A(n5375), .ZN(n3131) );
  NAND2_X1 U4300 ( .A1(n5570), .A2(n6607), .ZN(n5375) );
  OAI21_X1 U4301 ( .B1(n6096), .B2(n5570), .A(n5376), .ZN(n3130) );
  NAND2_X1 U4302 ( .A1(n5572), .A2(n6608), .ZN(n5376) );
  OAI21_X1 U4303 ( .B1(n6097), .B2(n5572), .A(n5377), .ZN(n3129) );
  NAND2_X1 U4304 ( .A1(n5570), .A2(n6609), .ZN(n5377) );
  OAI21_X1 U4305 ( .B1(n5525), .B2(n5572), .A(n5378), .ZN(n3128) );
  NAND2_X1 U4306 ( .A1(n5355), .A2(n6610), .ZN(n5378) );
  OAI21_X1 U4307 ( .B1(n6099), .B2(n5572), .A(n5379), .ZN(n3127) );
  NAND2_X1 U4308 ( .A1(n5355), .A2(n6611), .ZN(n5379) );
  OAI21_X1 U4309 ( .B1(n6100), .B2(n5572), .A(n5380), .ZN(n3126) );
  NAND2_X1 U4310 ( .A1(n5355), .A2(n6612), .ZN(n5380) );
  OAI21_X1 U4311 ( .B1(n6101), .B2(n5572), .A(n5381), .ZN(n3125) );
  NAND2_X1 U4312 ( .A1(n5355), .A2(n6613), .ZN(n5381) );
  OAI21_X1 U4313 ( .B1(n6102), .B2(n5572), .A(n5382), .ZN(n3124) );
  NAND2_X1 U4314 ( .A1(n5355), .A2(n6614), .ZN(n5382) );
  OAI21_X1 U4315 ( .B1(n6103), .B2(n5572), .A(n5383), .ZN(n3123) );
  NAND2_X1 U4316 ( .A1(n5355), .A2(n6615), .ZN(n5383) );
  OAI21_X1 U4317 ( .B1(n6104), .B2(n5572), .A(n5384), .ZN(n3122) );
  NAND2_X1 U4318 ( .A1(n5355), .A2(n6616), .ZN(n5384) );
  OAI21_X1 U4319 ( .B1(n6105), .B2(n5572), .A(n5385), .ZN(n3121) );
  NAND2_X1 U4320 ( .A1(n5355), .A2(n6617), .ZN(n5385) );
  OAI21_X1 U4321 ( .B1(n6106), .B2(n5572), .A(n5386), .ZN(n3120) );
  NAND2_X1 U4322 ( .A1(n5355), .A2(n6618), .ZN(n5386) );
  OAI21_X1 U4323 ( .B1(n6107), .B2(n5572), .A(n5387), .ZN(n3119) );
  NAND2_X1 U4324 ( .A1(n5355), .A2(n6619), .ZN(n5387) );
  NAND2_X1 U4325 ( .A1(n1777), .A2(n1521), .ZN(n5355) );
  NOR2_X1 U4326 ( .A1(n5388), .A2(n6066), .ZN(n1521) );
  OR2_X1 U4327 ( .A1(ADD_WR[1]), .A2(n6067), .ZN(n5388) );
  OAI21_X1 U4328 ( .B1(n6076), .B2(n5566), .A(n5390), .ZN(n3118) );
  NAND2_X1 U4329 ( .A1(n5566), .A2(n6516), .ZN(n5390) );
  OAI21_X1 U4330 ( .B1(n6077), .B2(n5562), .A(n5391), .ZN(n3117) );
  NAND2_X1 U4331 ( .A1(n5389), .A2(n6517), .ZN(n5391) );
  OAI21_X1 U4332 ( .B1(n6078), .B2(n5566), .A(n5392), .ZN(n3116) );
  NAND2_X1 U4333 ( .A1(n5562), .A2(n6518), .ZN(n5392) );
  OAI21_X1 U4334 ( .B1(n6079), .B2(n5562), .A(n5393), .ZN(n3115) );
  NAND2_X1 U4335 ( .A1(n5566), .A2(n6519), .ZN(n5393) );
  OAI21_X1 U4336 ( .B1(n6080), .B2(n5566), .A(n5394), .ZN(n3114) );
  NAND2_X1 U4337 ( .A1(n5562), .A2(n6520), .ZN(n5394) );
  OAI21_X1 U4338 ( .B1(n6081), .B2(n5562), .A(n5395), .ZN(n3113) );
  NAND2_X1 U4339 ( .A1(n5562), .A2(n6521), .ZN(n5395) );
  OAI21_X1 U4340 ( .B1(n5477), .B2(n5566), .A(n5396), .ZN(n3112) );
  NAND2_X1 U4341 ( .A1(n5562), .A2(n6522), .ZN(n5396) );
  OAI21_X1 U4342 ( .B1(n6083), .B2(n5562), .A(n5397), .ZN(n3111) );
  NAND2_X1 U4343 ( .A1(n5389), .A2(n6523), .ZN(n5397) );
  OAI21_X1 U4344 ( .B1(n6084), .B2(n5566), .A(n5398), .ZN(n3110) );
  NAND2_X1 U4345 ( .A1(n5389), .A2(n6524), .ZN(n5398) );
  OAI21_X1 U4346 ( .B1(n6085), .B2(n5562), .A(n5399), .ZN(n3109) );
  NAND2_X1 U4347 ( .A1(n5389), .A2(n6525), .ZN(n5399) );
  OAI21_X1 U4348 ( .B1(n6086), .B2(n5566), .A(n5400), .ZN(n3108) );
  NAND2_X1 U4349 ( .A1(n5389), .A2(n6526), .ZN(n5400) );
  OAI21_X1 U4350 ( .B1(n6087), .B2(n5566), .A(n5401), .ZN(n3107) );
  NAND2_X1 U4351 ( .A1(n5389), .A2(n6527), .ZN(n5401) );
  OAI21_X1 U4352 ( .B1(n6088), .B2(n5562), .A(n5402), .ZN(n3106) );
  NAND2_X1 U4353 ( .A1(n5389), .A2(n6528), .ZN(n5402) );
  OAI21_X1 U4354 ( .B1(n6089), .B2(n5562), .A(n5403), .ZN(n3105) );
  NAND2_X1 U4355 ( .A1(n5389), .A2(n6529), .ZN(n5403) );
  OAI21_X1 U4356 ( .B1(n6090), .B2(n5566), .A(n5404), .ZN(n3104) );
  NAND2_X1 U4357 ( .A1(n5389), .A2(n6530), .ZN(n5404) );
  OAI21_X1 U4358 ( .B1(n6091), .B2(n5562), .A(n5405), .ZN(n3103) );
  NAND2_X1 U4359 ( .A1(n5389), .A2(n6531), .ZN(n5405) );
  OAI21_X1 U4360 ( .B1(n5507), .B2(n5389), .A(n5406), .ZN(n3102) );
  NAND2_X1 U4361 ( .A1(n5562), .A2(n6532), .ZN(n5406) );
  OAI21_X1 U4362 ( .B1(n6093), .B2(n5389), .A(n5407), .ZN(n3101) );
  NAND2_X1 U4363 ( .A1(n5389), .A2(n6533), .ZN(n5407) );
  OAI21_X1 U4364 ( .B1(n6094), .B2(n5389), .A(n5408), .ZN(n3100) );
  NAND2_X1 U4365 ( .A1(n5562), .A2(n6534), .ZN(n5408) );
  OAI21_X1 U4366 ( .B1(n6095), .B2(n5389), .A(n5409), .ZN(n3099) );
  NAND2_X1 U4367 ( .A1(n5562), .A2(n6535), .ZN(n5409) );
  OAI21_X1 U4368 ( .B1(n6096), .B2(n5389), .A(n5410), .ZN(n3098) );
  NAND2_X1 U4369 ( .A1(n5562), .A2(n6536), .ZN(n5410) );
  OAI21_X1 U4370 ( .B1(n6097), .B2(n5389), .A(n5411), .ZN(n3097) );
  NAND2_X1 U4371 ( .A1(n5562), .A2(n6537), .ZN(n5411) );
  OAI21_X1 U4372 ( .B1(n5525), .B2(n5566), .A(n5412), .ZN(n3096) );
  NAND2_X1 U4373 ( .A1(n5562), .A2(n6538), .ZN(n5412) );
  OAI21_X1 U4374 ( .B1(n6099), .B2(n5566), .A(n5413), .ZN(n3095) );
  NAND2_X1 U4375 ( .A1(n5562), .A2(n6539), .ZN(n5413) );
  OAI21_X1 U4376 ( .B1(n6100), .B2(n5566), .A(n5414), .ZN(n3094) );
  NAND2_X1 U4377 ( .A1(n5562), .A2(n6540), .ZN(n5414) );
  OAI21_X1 U4378 ( .B1(n6101), .B2(n5566), .A(n5415), .ZN(n3093) );
  NAND2_X1 U4379 ( .A1(n5389), .A2(n6541), .ZN(n5415) );
  OAI21_X1 U4380 ( .B1(n6102), .B2(n5566), .A(n5416), .ZN(n3092) );
  NAND2_X1 U4381 ( .A1(n5389), .A2(n6542), .ZN(n5416) );
  OAI21_X1 U4382 ( .B1(n6103), .B2(n5566), .A(n5417), .ZN(n3091) );
  NAND2_X1 U4383 ( .A1(n5389), .A2(n6543), .ZN(n5417) );
  OAI21_X1 U4384 ( .B1(n6104), .B2(n5566), .A(n5418), .ZN(n3090) );
  NAND2_X1 U4385 ( .A1(n5389), .A2(n6544), .ZN(n5418) );
  OAI21_X1 U4386 ( .B1(n6105), .B2(n5566), .A(n5419), .ZN(n3089) );
  NAND2_X1 U4387 ( .A1(n5562), .A2(n6545), .ZN(n5419) );
  OAI21_X1 U4388 ( .B1(n6106), .B2(n5566), .A(n5420), .ZN(n3088) );
  NAND2_X1 U4389 ( .A1(n5389), .A2(n6546), .ZN(n5420) );
  OAI21_X1 U4390 ( .B1(n6107), .B2(n5389), .A(n5421), .ZN(n3087) );
  NAND2_X1 U4391 ( .A1(n5566), .A2(n6547), .ZN(n5421) );
  NAND2_X1 U4392 ( .A1(n2110), .A2(n1777), .ZN(n5389) );
  NOR2_X1 U4393 ( .A1(n5422), .A2(n6064), .ZN(n1777) );
  OR2_X1 U4394 ( .A1(n2273), .A2(n6065), .ZN(n5422) );
  NOR2_X1 U4395 ( .A1(n2453), .A2(ADD_WR[0]), .ZN(n2110) );
  OR2_X1 U4396 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .ZN(n2453) );
  OAI21_X1 U4397 ( .B1(n6076), .B2(n5558), .A(n5424), .ZN(n3086) );
  NAND2_X1 U4398 ( .A1(n5423), .A2(n6140), .ZN(n5424) );
  OAI21_X1 U4399 ( .B1(n6077), .B2(n5558), .A(n5425), .ZN(n3085) );
  NAND2_X1 U4400 ( .A1(n5423), .A2(n6141), .ZN(n5425) );
  OAI21_X1 U4401 ( .B1(n6078), .B2(n5558), .A(n5426), .ZN(n3084) );
  NAND2_X1 U4402 ( .A1(n5423), .A2(n6142), .ZN(n5426) );
  OAI21_X1 U4403 ( .B1(n6079), .B2(n5558), .A(n5427), .ZN(n3083) );
  NAND2_X1 U4404 ( .A1(n5423), .A2(n6143), .ZN(n5427) );
  OAI21_X1 U4405 ( .B1(n6080), .B2(n5558), .A(n5428), .ZN(n3082) );
  NAND2_X1 U4406 ( .A1(n5423), .A2(n6144), .ZN(n5428) );
  OAI21_X1 U4407 ( .B1(n6081), .B2(n5558), .A(n5429), .ZN(n3081) );
  NAND2_X1 U4408 ( .A1(n5423), .A2(n6145), .ZN(n5429) );
  OAI21_X1 U4409 ( .B1(n5477), .B2(n5558), .A(n5430), .ZN(n3080) );
  NAND2_X1 U4410 ( .A1(n5560), .A2(n6146), .ZN(n5430) );
  OAI21_X1 U4411 ( .B1(n6083), .B2(n5558), .A(n5431), .ZN(n3079) );
  NAND2_X1 U4412 ( .A1(n5558), .A2(n6147), .ZN(n5431) );
  OAI21_X1 U4413 ( .B1(n6084), .B2(n5558), .A(n5432), .ZN(n3078) );
  NAND2_X1 U4414 ( .A1(n5560), .A2(n6148), .ZN(n5432) );
  OAI21_X1 U4415 ( .B1(n6085), .B2(n5558), .A(n5433), .ZN(n3077) );
  NAND2_X1 U4416 ( .A1(n5558), .A2(n6149), .ZN(n5433) );
  OAI21_X1 U4417 ( .B1(n6086), .B2(n5558), .A(n5434), .ZN(n3076) );
  NAND2_X1 U4418 ( .A1(n5558), .A2(n6150), .ZN(n5434) );
  OAI21_X1 U4419 ( .B1(n6087), .B2(n5558), .A(n5435), .ZN(n3075) );
  NAND2_X1 U4420 ( .A1(n5423), .A2(n6151), .ZN(n5435) );
  OAI21_X1 U4421 ( .B1(n6088), .B2(n5560), .A(n5436), .ZN(n3074) );
  NAND2_X1 U4422 ( .A1(n5423), .A2(n6152), .ZN(n5436) );
  OAI21_X1 U4423 ( .B1(n6089), .B2(n5558), .A(n5437), .ZN(n3073) );
  NAND2_X1 U4424 ( .A1(n5423), .A2(n6153), .ZN(n5437) );
  OAI21_X1 U4425 ( .B1(n6090), .B2(n5560), .A(n5438), .ZN(n3072) );
  NAND2_X1 U4426 ( .A1(n5423), .A2(n6154), .ZN(n5438) );
  OAI21_X1 U4427 ( .B1(n6091), .B2(n5558), .A(n5439), .ZN(n3071) );
  NAND2_X1 U4428 ( .A1(n5423), .A2(n6155), .ZN(n5439) );
  OAI21_X1 U4429 ( .B1(n5507), .B2(n5560), .A(n5440), .ZN(n3070) );
  NAND2_X1 U4430 ( .A1(n5560), .A2(n6156), .ZN(n5440) );
  OAI21_X1 U4431 ( .B1(n6093), .B2(n5558), .A(n5441), .ZN(n3069) );
  NAND2_X1 U4432 ( .A1(n5423), .A2(n6157), .ZN(n5441) );
  OAI21_X1 U4433 ( .B1(n6094), .B2(n5560), .A(n5442), .ZN(n3068) );
  NAND2_X1 U4434 ( .A1(n5423), .A2(n6158), .ZN(n5442) );
  OAI21_X1 U4435 ( .B1(n6095), .B2(n5558), .A(n5443), .ZN(n3067) );
  NAND2_X1 U4436 ( .A1(n5558), .A2(n6159), .ZN(n5443) );
  OAI21_X1 U4437 ( .B1(n6096), .B2(n5560), .A(n5444), .ZN(n3066) );
  NAND2_X1 U4438 ( .A1(n5560), .A2(n6160), .ZN(n5444) );
  OAI21_X1 U4439 ( .B1(n6097), .B2(n5558), .A(n5445), .ZN(n3065) );
  NAND2_X1 U4440 ( .A1(n5560), .A2(n6161), .ZN(n5445) );
  OAI21_X1 U4441 ( .B1(n5525), .B2(n5560), .A(n5446), .ZN(n3064) );
  NAND2_X1 U4442 ( .A1(n5423), .A2(n6162), .ZN(n5446) );
  OAI21_X1 U4443 ( .B1(n6099), .B2(n5560), .A(n5447), .ZN(n3063) );
  NAND2_X1 U4444 ( .A1(n5423), .A2(n6163), .ZN(n5447) );
  OAI21_X1 U4445 ( .B1(n6100), .B2(n5560), .A(n5448), .ZN(n3062) );
  NAND2_X1 U4446 ( .A1(n5423), .A2(n6164), .ZN(n5448) );
  OAI21_X1 U4447 ( .B1(n6101), .B2(n5560), .A(n5449), .ZN(n3061) );
  NAND2_X1 U4448 ( .A1(n5423), .A2(n6165), .ZN(n5449) );
  OAI21_X1 U4449 ( .B1(n6102), .B2(n5560), .A(n5450), .ZN(n3060) );
  NAND2_X1 U4450 ( .A1(n5423), .A2(n6166), .ZN(n5450) );
  OAI21_X1 U4451 ( .B1(n6103), .B2(n5560), .A(n5451), .ZN(n3059) );
  NAND2_X1 U4452 ( .A1(n5423), .A2(n6167), .ZN(n5451) );
  OAI21_X1 U4453 ( .B1(n6104), .B2(n5560), .A(n5452), .ZN(n3058) );
  NAND2_X1 U4454 ( .A1(n5423), .A2(n6168), .ZN(n5452) );
  OAI21_X1 U4455 ( .B1(n6105), .B2(n5560), .A(n5453), .ZN(n3057) );
  NAND2_X1 U4456 ( .A1(n5423), .A2(n6169), .ZN(n5453) );
  OAI21_X1 U4457 ( .B1(n6106), .B2(n5560), .A(n5454), .ZN(n3056) );
  NAND2_X1 U4458 ( .A1(n5423), .A2(n6170), .ZN(n5454) );
  OAI21_X1 U4459 ( .B1(n6107), .B2(n5560), .A(n5455), .ZN(n3055) );
  NAND2_X1 U4460 ( .A1(n5423), .A2(n6171), .ZN(n5455) );
  NAND2_X1 U4461 ( .A1(n1812), .A2(n1520), .ZN(n5423) );
  NOR3_X1 U4462 ( .A1(n2273), .A2(ADD_WR[4]), .A3(ADD_WR[3]), .ZN(n1520) );
  NAND2_X1 U4463 ( .A1(WR), .A2(ENABLE), .ZN(n2273) );
  NOR2_X1 U4464 ( .A1(n5456), .A2(n6066), .ZN(n1812) );
  OR2_X1 U4465 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .ZN(n5456) );
  CLKBUF_X1 U2 ( .A(n5948), .Z(n6063) );
  CLKBUF_X1 U3 ( .A(n5948), .Z(n6062) );
  CLKBUF_X1 U6 ( .A(n5946), .Z(n6059) );
  CLKBUF_X1 U18 ( .A(n5949), .Z(n5948) );
  CLKBUF_X1 U20 ( .A(n5949), .Z(n5946) );
  CLKBUF_X1 U28 ( .A(n2148), .Z(n5807) );
  CLKBUF_X1 U44 ( .A(n2077), .Z(n5819) );
  CLKBUF_X1 U46 ( .A(n1846), .Z(n5861) );
  CLKBUF_X1 U50 ( .A(n1912), .Z(n5849) );
  CLKBUF_X1 U53 ( .A(n1744), .Z(n5880) );
  CLKBUF_X1 U54 ( .A(n1744), .Z(n5879) );
  CLKBUF_X1 U58 ( .A(n1487), .Z(n5928) );
  CLKBUF_X1 U59 ( .A(n1487), .Z(n5929) );
  CLKBUF_X1 U60 ( .A(n2148), .Z(n5809) );
  CLKBUF_X1 U67 ( .A(n2077), .Z(n5821) );
  CLKBUF_X1 U68 ( .A(n1846), .Z(n5863) );
  CLKBUF_X1 U70 ( .A(n1912), .Z(n5851) );
  CLKBUF_X1 U76 ( .A(n1591), .Z(n5910) );
  CLKBUF_X1 U81 ( .A(n2308), .Z(n5783) );
  CLKBUF_X1 U88 ( .A(n5389), .Z(n5562) );
  CLKBUF_X1 U98 ( .A(n1828), .Z(n5868) );
  CLKBUF_X1 U100 ( .A(n1659), .Z(n5898) );
  CLKBUF_X1 U106 ( .A(n2308), .Z(n5785) );
  CLKBUF_X1 U121 ( .A(n1779), .Z(n5877) );
  CLKBUF_X1 U122 ( .A(n1779), .Z(n5876) );
  CLKBUF_X1 U126 ( .A(n2011), .Z(n5835) );
  CLKBUF_X1 U128 ( .A(n2044), .Z(n5829) );
  CLKBUF_X1 U131 ( .A(n1625), .Z(n5907) );
  CLKBUF_X1 U132 ( .A(n1625), .Z(n5906) );
  CLKBUF_X1 U138 ( .A(n1557), .Z(n5918) );
  CLKBUF_X1 U140 ( .A(n1522), .Z(n5924) );
  CLKBUF_X1 U142 ( .A(n2189), .Z(n5805) );
  CLKBUF_X1 U144 ( .A(n2231), .Z(n5799) );
  CLKBUF_X1 U146 ( .A(n2274), .Z(n5793) );
  CLKBUF_X1 U150 ( .A(n5423), .Z(n5558) );
  CLKBUF_X1 U152 ( .A(n2342), .Z(n5781) );
  CLKBUF_X1 U154 ( .A(n2386), .Z(n5775) );
  CLKBUF_X1 U156 ( .A(n2420), .Z(n5769) );
  CLKBUF_X1 U160 ( .A(n1879), .Z(n5859) );
  CLKBUF_X1 U162 ( .A(n5355), .Z(n5570) );
  CLKBUF_X1 U165 ( .A(n1945), .Z(n5846) );
  CLKBUF_X1 U166 ( .A(n1945), .Z(n5847) );
  CLKBUF_X1 U170 ( .A(n1693), .Z(n5894) );
  CLKBUF_X1 U171 ( .A(n1726), .Z(n5889) );
  CLKBUF_X1 U172 ( .A(n1726), .Z(n5888) );
  CLKBUF_X1 U173 ( .A(n1978), .Z(n5840) );
  CLKBUF_X1 U174 ( .A(n1978), .Z(n5841) );
  CLKBUF_X1 U180 ( .A(n2111), .Z(n5817) );
  CLKBUF_X1 U182 ( .A(n2274), .Z(n5794) );
  CLKBUF_X1 U184 ( .A(n5423), .Z(n5560) );
  CLKBUF_X1 U185 ( .A(n2342), .Z(n5782) );
  CLKBUF_X1 U186 ( .A(n2386), .Z(n5776) );
  CLKBUF_X1 U187 ( .A(n2420), .Z(n5770) );
  CLKBUF_X1 U189 ( .A(n5389), .Z(n5566) );
  CLKBUF_X1 U190 ( .A(n2011), .Z(n5836) );
  CLKBUF_X1 U191 ( .A(n2044), .Z(n5830) );
  CLKBUF_X1 U194 ( .A(n1591), .Z(n5914) );
  CLKBUF_X1 U196 ( .A(n1557), .Z(n5920) );
  CLKBUF_X1 U197 ( .A(n1522), .Z(n5926) );
  CLKBUF_X1 U198 ( .A(n2189), .Z(n5806) );
  CLKBUF_X1 U199 ( .A(n2231), .Z(n5800) );
  CLKBUF_X1 U201 ( .A(n1879), .Z(n5860) );
  CLKBUF_X1 U202 ( .A(n5355), .Z(n5572) );
  CLKBUF_X1 U206 ( .A(n1693), .Z(n5896) );
  CLKBUF_X1 U209 ( .A(n1828), .Z(n5872) );
  CLKBUF_X1 U210 ( .A(n1659), .Z(n5902) );
  CLKBUF_X1 U211 ( .A(n2111), .Z(n5818) );
  CLKBUF_X1 U212 ( .A(n5458), .Z(n5457) );
  CLKBUF_X1 U213 ( .A(n5939), .Z(n5458) );
  CLKBUF_X1 U214 ( .A(RESET), .Z(n5949) );
  INV_X1 U219 ( .A(ENABLE), .ZN(n5939) );
  CLKBUF_X1 U226 ( .A(n4461), .Z(n5634) );
  CLKBUF_X1 U230 ( .A(n2477), .Z(n5735) );
  CLKBUF_X1 U246 ( .A(n4453), .Z(n5645) );
  CLKBUF_X1 U257 ( .A(n2502), .Z(n5691) );
  CLKBUF_X1 U278 ( .A(n2483), .Z(n5717) );
  CLKBUF_X1 U283 ( .A(n4444), .Z(n5664) );
  CLKBUF_X1 U302 ( .A(n4485), .Z(n5591) );
  CLKBUF_X1 U305 ( .A(n4493), .Z(n5573) );
  CLKBUF_X1 U321 ( .A(n2505), .Z(n5681) );
  CLKBUF_X1 U329 ( .A(n2492), .Z(n5709) );
  CLKBUF_X1 U337 ( .A(n4481), .Z(n5598) );
  CLKBUF_X1 U349 ( .A(n2460), .Z(n5763) );
  CLKBUF_X1 U351 ( .A(n4447), .Z(n5659) );
  CLKBUF_X1 U352 ( .A(n4486), .Z(n5590) );
  CLKBUF_X1 U353 ( .A(n4492), .Z(n5578) );
  CLKBUF_X1 U355 ( .A(n2479), .Z(n5731) );
  CLKBUF_X1 U356 ( .A(n2465), .Z(n5755) );
  CLKBUF_X1 U357 ( .A(n2493), .Z(n5707) );
  CLKBUF_X1 U358 ( .A(n2504), .Z(n5686) );
  CLKBUF_X1 U359 ( .A(n2510), .Z(n5674) );
  CLKBUF_X1 U360 ( .A(n4480), .Z(n5602) );
  CLKBUF_X1 U361 ( .A(n2498), .Z(n5698) );
  CLKBUF_X1 U363 ( .A(n4451), .Z(n5653) );
  CLKBUF_X1 U364 ( .A(n4484), .Z(n5596) );
  CLKBUF_X1 U365 ( .A(n2471), .Z(n5743) );
  CLKBUF_X1 U366 ( .A(n2469), .Z(n5749) );
  CLKBUF_X1 U368 ( .A(n4463), .Z(n5629) );
  CLKBUF_X1 U369 ( .A(n4473), .Z(n5617) );
  CLKBUF_X1 U370 ( .A(n4475), .Z(n5611) );
  CLKBUF_X1 U371 ( .A(n4490), .Z(n5584) );
  CLKBUF_X1 U372 ( .A(n2481), .Z(n5725) );
  CLKBUF_X1 U373 ( .A(n2491), .Z(n5713) );
  CLKBUF_X1 U374 ( .A(n2508), .Z(n5680) );
  CLKBUF_X1 U375 ( .A(n4459), .Z(n5641) );
  CLKBUF_X1 U376 ( .A(n4465), .Z(n5623) );
  CLKBUF_X1 U377 ( .A(n4478), .Z(n5608) );
  CLKBUF_X1 U379 ( .A(n2496), .Z(n5704) );
  CLKBUF_X1 U381 ( .A(n2462), .Z(n5761) );
  CLKBUF_X1 U382 ( .A(n4462), .Z(n5632) );
  CLKBUF_X1 U383 ( .A(n4454), .Z(n5644) );
  CLKBUF_X1 U384 ( .A(n4479), .Z(n5605) );
  CLKBUF_X1 U385 ( .A(n2480), .Z(n5728) );
  CLKBUF_X1 U386 ( .A(n2497), .Z(n5701) );
  CLKBUF_X1 U387 ( .A(n4464), .Z(n5626) );
  CLKBUF_X1 U388 ( .A(n4448), .Z(n5656) );
  CLKBUF_X1 U389 ( .A(n4474), .Z(n5614) );
  CLKBUF_X1 U391 ( .A(n4487), .Z(n5587) );
  CLKBUF_X1 U392 ( .A(n2466), .Z(n5752) );
  CLKBUF_X1 U393 ( .A(n2472), .Z(n5740) );
  CLKBUF_X1 U395 ( .A(n2503), .Z(n5689) );
  CLKBUF_X1 U397 ( .A(n4460), .Z(n5638) );
  CLKBUF_X1 U398 ( .A(n4466), .Z(n5620) );
  CLKBUF_X1 U399 ( .A(n4491), .Z(n5581) );
  CLKBUF_X1 U401 ( .A(n2478), .Z(n5734) );
  CLKBUF_X1 U402 ( .A(n2482), .Z(n5722) );
  CLKBUF_X1 U403 ( .A(n2484), .Z(n5716) );
  CLKBUF_X1 U404 ( .A(n2509), .Z(n5677) );
  CLKBUF_X1 U405 ( .A(n2511), .Z(n5671) );
  CLKBUF_X1 U406 ( .A(n4452), .Z(n5650) );
  CLKBUF_X1 U408 ( .A(n2470), .Z(n5746) );
  CLKBUF_X1 U409 ( .A(n2499), .Z(n5695) );
  CLKBUF_X1 U410 ( .A(n4445), .Z(n5662) );
  CLKBUF_X1 U411 ( .A(n2463), .Z(n5758) );
  CLKBUF_X1 U412 ( .A(n4442), .Z(n5668) );
  CLKBUF_X1 U429 ( .A(n6077), .Z(n5463) );
  CLKBUF_X1 U433 ( .A(n6105), .Z(n5547) );
  CLKBUF_X1 U445 ( .A(n6093), .Z(n5511) );
  CLKBUF_X1 U455 ( .A(n6098), .Z(n5525) );
  CLKBUF_X1 U461 ( .A(n6092), .Z(n5507) );
  CLKBUF_X1 U471 ( .A(n6082), .Z(n5477) );
  CLKBUF_X1 U478 ( .A(n6107), .Z(n5554) );
  CLKBUF_X1 U479 ( .A(n6106), .Z(n5551) );
  CLKBUF_X1 U481 ( .A(n6104), .Z(n5545) );
  CLKBUF_X1 U482 ( .A(n6103), .Z(n5542) );
  CLKBUF_X1 U483 ( .A(n6102), .Z(n5539) );
  CLKBUF_X1 U484 ( .A(n6101), .Z(n5536) );
  CLKBUF_X1 U485 ( .A(n6100), .Z(n5533) );
  CLKBUF_X1 U486 ( .A(n6099), .Z(n5530) );
  CLKBUF_X1 U488 ( .A(n6097), .Z(n5524) );
  CLKBUF_X1 U489 ( .A(n6096), .Z(n5521) );
  CLKBUF_X1 U490 ( .A(n6095), .Z(n5518) );
  CLKBUF_X1 U491 ( .A(n6094), .Z(n5515) );
  CLKBUF_X1 U494 ( .A(n6091), .Z(n5506) );
  CLKBUF_X1 U495 ( .A(n6090), .Z(n5503) );
  CLKBUF_X1 U496 ( .A(n6089), .Z(n5500) );
  CLKBUF_X1 U497 ( .A(n6088), .Z(n5497) );
  CLKBUF_X1 U498 ( .A(n6087), .Z(n5494) );
  CLKBUF_X1 U499 ( .A(n6086), .Z(n5491) );
  CLKBUF_X1 U500 ( .A(n6085), .Z(n5488) );
  CLKBUF_X1 U501 ( .A(n6084), .Z(n5485) );
  CLKBUF_X1 U502 ( .A(n6083), .Z(n5482) );
  CLKBUF_X1 U504 ( .A(n6081), .Z(n5476) );
  CLKBUF_X1 U505 ( .A(n6080), .Z(n5473) );
  CLKBUF_X1 U506 ( .A(n6079), .Z(n5470) );
  CLKBUF_X1 U507 ( .A(n6078), .Z(n5467) );
  CLKBUF_X1 U509 ( .A(n6076), .Z(n5461) );
  INV_X1 U511 ( .A(ADD_WR[0]), .ZN(n6067) );
  INV_X1 U512 ( .A(ADD_WR[2]), .ZN(n6066) );
  INV_X1 U514 ( .A(ADD_WR[4]), .ZN(n6064) );
  INV_X1 U515 ( .A(ADD_WR[3]), .ZN(n6065) );
  INV_X1 U516 ( .A(DATAIN[10]), .ZN(n6097) );
  INV_X1 U517 ( .A(DATAIN[11]), .ZN(n6096) );
  INV_X1 U518 ( .A(DATAIN[12]), .ZN(n6095) );
  INV_X1 U519 ( .A(DATAIN[13]), .ZN(n6094) );
  INV_X1 U520 ( .A(DATAIN[14]), .ZN(n6093) );
  INV_X1 U521 ( .A(DATAIN[8]), .ZN(n6099) );
  INV_X1 U522 ( .A(DATAIN[9]), .ZN(n6098) );
  INV_X1 U523 ( .A(DATAIN[30]), .ZN(n6077) );
  INV_X1 U524 ( .A(DATAIN[31]), .ZN(n6076) );
  INV_X1 U557 ( .A(ADD_RD2[0]), .ZN(n6075) );
  INV_X1 U558 ( .A(ADD_RD1[0]), .ZN(n6071) );
  INV_X1 U559 ( .A(WR), .ZN(n6620) );
  INV_X1 U4466 ( .A(ADD_RD2[4]), .ZN(n6072) );
  INV_X1 U4467 ( .A(ADD_RD1[4]), .ZN(n6068) );
  INV_X1 U4948 ( .A(DATAIN[0]), .ZN(n6107) );
  INV_X1 U4949 ( .A(DATAIN[1]), .ZN(n6106) );
  INV_X1 U4950 ( .A(DATAIN[15]), .ZN(n6092) );
  INV_X1 U4951 ( .A(DATAIN[16]), .ZN(n6091) );
  INV_X1 U4952 ( .A(DATAIN[17]), .ZN(n6090) );
  INV_X1 U4953 ( .A(DATAIN[18]), .ZN(n6089) );
  INV_X1 U4954 ( .A(DATAIN[19]), .ZN(n6088) );
  INV_X1 U4955 ( .A(DATAIN[20]), .ZN(n6087) );
  INV_X1 U4956 ( .A(DATAIN[21]), .ZN(n6086) );
  INV_X1 U4957 ( .A(DATAIN[22]), .ZN(n6085) );
  INV_X1 U4958 ( .A(DATAIN[23]), .ZN(n6084) );
  INV_X1 U4959 ( .A(DATAIN[24]), .ZN(n6083) );
  INV_X1 U4960 ( .A(DATAIN[25]), .ZN(n6082) );
  INV_X1 U4961 ( .A(DATAIN[26]), .ZN(n6081) );
  INV_X1 U4962 ( .A(DATAIN[27]), .ZN(n6080) );
  INV_X1 U4963 ( .A(DATAIN[28]), .ZN(n6079) );
  INV_X1 U4964 ( .A(DATAIN[29]), .ZN(n6078) );
  INV_X1 U4965 ( .A(DATAIN[2]), .ZN(n6105) );
  INV_X1 U4966 ( .A(DATAIN[3]), .ZN(n6104) );
  INV_X1 U4967 ( .A(DATAIN[4]), .ZN(n6103) );
  INV_X1 U4968 ( .A(DATAIN[5]), .ZN(n6102) );
  INV_X1 U4969 ( .A(DATAIN[6]), .ZN(n6101) );
  INV_X1 U4970 ( .A(DATAIN[7]), .ZN(n6100) );
  INV_X1 U4971 ( .A(ADD_RD2[2]), .ZN(n6073) );
  INV_X1 U4972 ( .A(ADD_RD2[1]), .ZN(n6074) );
  INV_X1 U4973 ( .A(ADD_RD1[2]), .ZN(n6069) );
  INV_X1 U4974 ( .A(ADD_RD1[1]), .ZN(n6070) );
  CLKBUF_X1 U4976 ( .A(n6063), .Z(n5952) );
  CLKBUF_X1 U4977 ( .A(n6063), .Z(n5953) );
  CLKBUF_X1 U4978 ( .A(n6063), .Z(n5954) );
  CLKBUF_X1 U4979 ( .A(n6063), .Z(n5955) );
  CLKBUF_X1 U4980 ( .A(n6063), .Z(n5956) );
  CLKBUF_X1 U4981 ( .A(n6063), .Z(n5957) );
  CLKBUF_X1 U4982 ( .A(n6062), .Z(n5958) );
  CLKBUF_X1 U4983 ( .A(n6062), .Z(n5959) );
  CLKBUF_X1 U4984 ( .A(n6062), .Z(n5960) );
  CLKBUF_X1 U4985 ( .A(n6062), .Z(n5961) );
  CLKBUF_X1 U4986 ( .A(n6062), .Z(n5962) );
  CLKBUF_X1 U4987 ( .A(n6062), .Z(n5963) );
  CLKBUF_X1 U4998 ( .A(n5949), .Z(n5974) );
  CLKBUF_X1 U5006 ( .A(n6063), .Z(n5982) );
  CLKBUF_X1 U5007 ( .A(n5949), .Z(n5983) );
  CLKBUF_X1 U5008 ( .A(n5946), .Z(n5984) );
  CLKBUF_X1 U5009 ( .A(n6059), .Z(n5985) );
  CLKBUF_X1 U5016 ( .A(n6063), .Z(n5992) );
  CLKBUF_X1 U5017 ( .A(n6062), .Z(n5993) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n3230), .CK(CLK), .RN(n5955), .Q(n640)
         );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n3231), .CK(CLK), .RN(n5956), .Q(n639)
         );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n3232), .CK(CLK), .RN(n5957), .Q(n638)
         );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n3233), .CK(CLK), .RN(n5958), .Q(n637)
         );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n3234), .CK(CLK), .RN(n5959), .Q(n636)
         );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n3235), .CK(CLK), .RN(n5960), .Q(n635)
         );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n3236), .CK(CLK), .RN(n5961), .Q(n634)
         );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n3237), .CK(CLK), .RN(n5962), .Q(n633)
         );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n3238), .CK(CLK), .RN(n5963), .Q(n632)
         );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n3239), .CK(CLK), .RN(RESET), .Q(n631)
         );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n3240), .CK(CLK), .RN(RESET), .Q(n630)
         );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n3241), .CK(CLK), .RN(RESET), .Q(n629)
         );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n3242), .CK(CLK), .RN(RESET), .Q(n628)
         );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n3243), .CK(CLK), .RN(RESET), .Q(n627)
         );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n3244), .CK(CLK), .RN(RESET), .Q(n626)
         );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n3245), .CK(CLK), .RN(RESET), .Q(n625)
         );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n3246), .CK(CLK), .RN(RESET), .Q(n624)
         );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n3247), .CK(CLK), .RN(RESET), .Q(n623)
         );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n3248), .CK(CLK), .RN(RESET), .Q(n622)
         );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n3249), .CK(CLK), .RN(n5974), .Q(n621)
         );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n3250), .CK(CLK), .RN(RESET), .Q(n620)
         );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n3251), .CK(CLK), .RN(RESET), .Q(n619)
         );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n3252), .CK(CLK), .RN(RESET), .Q(n618) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n3253), .CK(CLK), .RN(RESET), .Q(n617) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n3254), .CK(CLK), .RN(RESET), .Q(n616) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3255), .CK(CLK), .RN(RESET), .Q(n615) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3256), .CK(CLK), .RN(RESET), .Q(n614) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3257), .CK(CLK), .RN(n5982), .Q(n613) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3258), .CK(CLK), .RN(n5983), .Q(n612) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n3259), .CK(CLK), .RN(n5984), .Q(n611) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n3260), .CK(CLK), .RN(n5985), .Q(n610) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3261), .CK(CLK), .RN(RESET), .Q(n609) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3262), .CK(CLK), .RN(RESET), .Q(n6108)
         );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3263), .CK(CLK), .RN(n5948), .Q(n6109)
         );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3264), .CK(CLK), .RN(n5953), .Q(n6110)
         );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3265), .CK(CLK), .RN(n5992), .Q(n6111)
         );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3266), .CK(CLK), .RN(n5958), .Q(n6112)
         );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3267), .CK(CLK), .RN(RESET), .Q(n6113)
         );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3268), .CK(CLK), .RN(n5949), .Q(n6114)
         );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3269), .CK(CLK), .RN(n5948), .Q(n6115)
         );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3270), .CK(CLK), .RN(RESET), .Q(n6116)
         );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3271), .CK(CLK), .RN(RESET), .Q(n6117)
         );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3272), .CK(CLK), .RN(n5953), .Q(n6118)
         );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3273), .CK(CLK), .RN(n5957), .Q(n6119)
         );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3274), .CK(CLK), .RN(n5992), .Q(n6120)
         );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3275), .CK(CLK), .RN(n5982), .Q(n6121)
         );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3276), .CK(CLK), .RN(n6062), .Q(n6122)
         );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3277), .CK(CLK), .RN(RESET), .Q(n6123)
         );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3278), .CK(CLK), .RN(n6059), .Q(n6124)
         );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3279), .CK(CLK), .RN(RESET), .Q(n6125)
         );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3280), .CK(CLK), .RN(RESET), .Q(n6126)
         );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3281), .CK(CLK), .RN(n6062), .Q(n6127)
         );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3282), .CK(CLK), .RN(n5957), .Q(n6128)
         );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3283), .CK(CLK), .RN(n6059), .Q(n6129)
         );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3284), .CK(CLK), .RN(n6063), .Q(n6130)
         );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3285), .CK(CLK), .RN(RESET), .Q(n6131)
         );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3286), .CK(CLK), .RN(n5946), .Q(n6132)
         );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3287), .CK(CLK), .RN(n5954), .Q(n6133)
         );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3288), .CK(CLK), .RN(n6062), .Q(n6134)
         );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3289), .CK(CLK), .RN(n5948), .Q(n6135)
         );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3290), .CK(CLK), .RN(RESET), .Q(n6136)
         );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3291), .CK(CLK), .RN(n5946), .Q(n6137)
         );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3292), .CK(CLK), .RN(n6062), .Q(n6138)
         );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3293), .CK(CLK), .RN(n5948), .Q(n6139)
         );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3294), .CK(CLK), .RN(RESET), .Q(n608)
         );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3295), .CK(CLK), .RN(n5946), .Q(n607)
         );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3296), .CK(CLK), .RN(n5984), .Q(n606)
         );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3297), .CK(CLK), .RN(n5949), .Q(n605)
         );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3298), .CK(CLK), .RN(n6062), .Q(n604)
         );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3299), .CK(CLK), .RN(n5985), .Q(n603)
         );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3300), .CK(CLK), .RN(n5949), .Q(n602)
         );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3301), .CK(CLK), .RN(n5957), .Q(n601)
         );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3302), .CK(CLK), .RN(n5949), .Q(n600)
         );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3303), .CK(CLK), .RN(n5949), .Q(n599)
         );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3304), .CK(CLK), .RN(n5949), .Q(n598)
         );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3305), .CK(CLK), .RN(n5949), .Q(n597)
         );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3306), .CK(CLK), .RN(n5949), .Q(n596)
         );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3307), .CK(CLK), .RN(RESET), .Q(n595)
         );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3308), .CK(CLK), .RN(n5953), .Q(n594)
         );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3309), .CK(CLK), .RN(RESET), .Q(n593)
         );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3310), .CK(CLK), .RN(RESET), .Q(n592)
         );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3311), .CK(CLK), .RN(n5982), .Q(n591)
         );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3312), .CK(CLK), .RN(n5983), .Q(n590)
         );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3313), .CK(CLK), .RN(n5984), .Q(n589)
         );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3314), .CK(CLK), .RN(n5985), .Q(n588)
         );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3315), .CK(CLK), .RN(RESET), .Q(n587)
         );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3316), .CK(CLK), .RN(RESET), .Q(n586) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3317), .CK(CLK), .RN(n5953), .Q(n585) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3318), .CK(CLK), .RN(RESET), .Q(n584) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3319), .CK(CLK), .RN(n5993), .Q(n583) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3320), .CK(CLK), .RN(RESET), .Q(n582) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3321), .CK(CLK), .RN(n5954), .Q(n581) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3322), .CK(CLK), .RN(n5982), .Q(n580) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3323), .CK(CLK), .RN(n5955), .Q(n579) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3324), .CK(CLK), .RN(n5983), .Q(n578) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3325), .CK(CLK), .RN(n5956), .Q(n577) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n3086), .CK(CLK), .RN(n5984), .Q(n6140)
         );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n3085), .CK(CLK), .RN(n5985), .Q(n6141)
         );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n3084), .CK(CLK), .RN(RESET), .Q(n6142)
         );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n3083), .CK(CLK), .RN(RESET), .Q(n6143)
         );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n3082), .CK(CLK), .RN(RESET), .Q(n6144)
         );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n3081), .CK(CLK), .RN(n5993), .Q(n6145)
         );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n3080), .CK(CLK), .RN(n5974), .Q(n6146)
         );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n3079), .CK(CLK), .RN(n5952), .Q(n6147)
         );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n3078), .CK(CLK), .RN(RESET), .Q(n6148)
         );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n3077), .CK(CLK), .RN(RESET), .Q(n6149)
         );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n3076), .CK(CLK), .RN(n5949), .Q(n6150)
         );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n3075), .CK(CLK), .RN(RESET), .Q(n6151)
         );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n3074), .CK(CLK), .RN(RESET), .Q(n6152)
         );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n3073), .CK(CLK), .RN(RESET), .Q(n6153)
         );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n3072), .CK(CLK), .RN(RESET), .Q(n6154)
         );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n3071), .CK(CLK), .RN(RESET), .Q(n6155)
         );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n3070), .CK(CLK), .RN(n6059), .Q(n6156)
         );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n3069), .CK(CLK), .RN(RESET), .Q(n6157)
         );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n3068), .CK(CLK), .RN(n6059), .Q(n6158)
         );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n3067), .CK(CLK), .RN(n5956), .Q(n6159)
         );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n3066), .CK(CLK), .RN(n5985), .Q(n6160)
         );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n3065), .CK(CLK), .RN(n5948), .Q(n6161)
         );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n3064), .CK(CLK), .RN(n5952), .Q(n6162)
         );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n3063), .CK(CLK), .RN(n5959), .Q(n6163)
         );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n3062), .CK(CLK), .RN(RESET), .Q(n6164)
         );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n3061), .CK(CLK), .RN(n5983), .Q(n6165)
         );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n3060), .CK(CLK), .RN(n5952), .Q(n6166)
         );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n3059), .CK(CLK), .RN(n6063), .Q(n6167)
         );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n3058), .CK(CLK), .RN(n6059), .Q(n6168)
         );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n3057), .CK(CLK), .RN(RESET), .Q(n6169)
         );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n3056), .CK(CLK), .RN(RESET), .Q(n6170)
         );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n3055), .CK(CLK), .RN(n6062), .Q(n6171)
         );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n4189), .CK(CLK), .RN(n5946), .Q(n6172)
         );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n4188), .CK(CLK), .RN(RESET), .Q(n6173)
         );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n4187), .CK(CLK), .RN(n5958), .Q(n6174)
         );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n4186), .CK(CLK), .RN(n5982), .Q(n6175)
         );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n4185), .CK(CLK), .RN(n5957), .Q(n6176)
         );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n4184), .CK(CLK), .RN(n5946), .Q(n6177)
         );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n4183), .CK(CLK), .RN(n5957), .Q(n6178)
         );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n4182), .CK(CLK), .RN(n5992), .Q(n6179)
         );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n4181), .CK(CLK), .RN(n5993), .Q(n6180)
         );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n4180), .CK(CLK), .RN(RESET), .Q(n6181)
         );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n4179), .CK(CLK), .RN(RESET), .Q(n6182)
         );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n4178), .CK(CLK), .RN(RESET), .Q(n6183)
         );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n4177), .CK(CLK), .RN(n5974), .Q(n6184)
         );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n4176), .CK(CLK), .RN(RESET), .Q(n6185)
         );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n4175), .CK(CLK), .RN(n5955), .Q(n6186)
         );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n4174), .CK(CLK), .RN(n6063), .Q(n6187)
         );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n4173), .CK(CLK), .RN(n5949), .Q(n6188)
         );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n4172), .CK(CLK), .RN(RESET), .Q(n6189)
         );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n4171), .CK(CLK), .RN(RESET), .Q(n6190)
         );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n4170), .CK(CLK), .RN(n5992), .Q(n6191)
         );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n4169), .CK(CLK), .RN(RESET), .Q(n6192)
         );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n4168), .CK(CLK), .RN(n5956), .Q(n6193)
         );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n4167), .CK(CLK), .RN(n6059), .Q(n6194)
         );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n4166), .CK(CLK), .RN(RESET), .Q(n6195)
         );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n4165), .CK(CLK), .RN(n5985), .Q(n6196)
         );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n4164), .CK(CLK), .RN(n5956), .Q(n6197)
         );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n4163), .CK(CLK), .RN(RESET), .Q(n6198)
         );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n4162), .CK(CLK), .RN(n5959), .Q(n6199)
         );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n4161), .CK(CLK), .RN(n5949), .Q(n6200)
         );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n4160), .CK(CLK), .RN(RESET), .Q(n6201)
         );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n4159), .CK(CLK), .RN(n5949), .Q(n6202)
         );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n4158), .CK(CLK), .RN(n5961), .Q(n6203)
         );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3326), .CK(CLK), .RN(n5949), .Q(n6204)
         );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3327), .CK(CLK), .RN(n5953), .Q(n6205)
         );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3328), .CK(CLK), .RN(n5949), .Q(n6206)
         );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3329), .CK(CLK), .RN(n5960), .Q(n6207)
         );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3330), .CK(CLK), .RN(RESET), .Q(n6208)
         );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3331), .CK(CLK), .RN(RESET), .Q(n6209)
         );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3332), .CK(CLK), .RN(n5953), .Q(n6210)
         );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3333), .CK(CLK), .RN(RESET), .Q(n6211)
         );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3334), .CK(CLK), .RN(RESET), .Q(n6212)
         );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3335), .CK(CLK), .RN(n5953), .Q(n6213)
         );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3336), .CK(CLK), .RN(n5953), .Q(n6214)
         );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3337), .CK(CLK), .RN(RESET), .Q(n6215)
         );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3338), .CK(CLK), .RN(RESET), .Q(n6216)
         );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3339), .CK(CLK), .RN(n5953), .Q(n6217)
         );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3340), .CK(CLK), .RN(RESET), .Q(n6218)
         );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3341), .CK(CLK), .RN(RESET), .Q(n6219)
         );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3342), .CK(CLK), .RN(RESET), .Q(n6220)
         );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3343), .CK(CLK), .RN(n5953), .Q(n6221)
         );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3344), .CK(CLK), .RN(RESET), .Q(n6222)
         );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3345), .CK(CLK), .RN(RESET), .Q(n6223)
         );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3346), .CK(CLK), .RN(RESET), .Q(n6224)
         );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3347), .CK(CLK), .RN(n5953), .Q(n6225)
         );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3348), .CK(CLK), .RN(RESET), .Q(n6226)
         );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3349), .CK(CLK), .RN(RESET), .Q(n6227)
         );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3350), .CK(CLK), .RN(n5953), .Q(n6228)
         );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3351), .CK(CLK), .RN(RESET), .Q(n6229)
         );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3352), .CK(CLK), .RN(RESET), .Q(n6230)
         );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3353), .CK(CLK), .RN(RESET), .Q(n6231)
         );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3354), .CK(CLK), .RN(n5982), .Q(n6232)
         );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3355), .CK(CLK), .RN(n5983), .Q(n6233)
         );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3356), .CK(CLK), .RN(n5984), .Q(n6234)
         );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3357), .CK(CLK), .RN(n5985), .Q(n6235)
         );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3358), .CK(CLK), .RN(RESET), .Q(n480)
         );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3359), .CK(CLK), .RN(RESET), .Q(n479)
         );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3360), .CK(CLK), .RN(n6063), .Q(n478)
         );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3361), .CK(CLK), .RN(n5952), .Q(n477)
         );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3362), .CK(CLK), .RN(n5954), .Q(n476)
         );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3363), .CK(CLK), .RN(n5955), .Q(n475)
         );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3364), .CK(CLK), .RN(n5959), .Q(n474)
         );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3365), .CK(CLK), .RN(n5960), .Q(n473)
         );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3366), .CK(CLK), .RN(n5961), .Q(n472)
         );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3367), .CK(CLK), .RN(n5962), .Q(n471)
         );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3368), .CK(CLK), .RN(n5963), .Q(n470)
         );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3369), .CK(CLK), .RN(RESET), .Q(n469)
         );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3370), .CK(CLK), .RN(RESET), .Q(n468)
         );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3371), .CK(CLK), .RN(RESET), .Q(n467)
         );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3372), .CK(CLK), .RN(RESET), .Q(n466)
         );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3373), .CK(CLK), .RN(RESET), .Q(n465)
         );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3374), .CK(CLK), .RN(RESET), .Q(n464)
         );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3375), .CK(CLK), .RN(n5958), .Q(n463)
         );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3376), .CK(CLK), .RN(n6062), .Q(n462)
         );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3377), .CK(CLK), .RN(n6059), .Q(n461)
         );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3378), .CK(CLK), .RN(RESET), .Q(n460)
         );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3379), .CK(CLK), .RN(RESET), .Q(n459)
         );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3380), .CK(CLK), .RN(RESET), .Q(n458) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3381), .CK(CLK), .RN(RESET), .Q(n457) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3382), .CK(CLK), .RN(n5974), .Q(n456) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3383), .CK(CLK), .RN(RESET), .Q(n455) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3384), .CK(CLK), .RN(RESET), .Q(n454) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3385), .CK(CLK), .RN(RESET), .Q(n453) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3386), .CK(CLK), .RN(n5993), .Q(n452) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3387), .CK(CLK), .RN(n6063), .Q(n451) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3388), .CK(CLK), .RN(RESET), .Q(n450) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3389), .CK(CLK), .RN(n5954), .Q(n449) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n3390), .CK(CLK), .RN(RESET), .Q(n576)
         );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n3391), .CK(CLK), .RN(RESET), .Q(n575)
         );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n3392), .CK(CLK), .RN(n5956), .Q(n574)
         );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n3393), .CK(CLK), .RN(n5993), .Q(n573)
         );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n3394), .CK(CLK), .RN(RESET), .Q(n572)
         );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n3395), .CK(CLK), .RN(RESET), .Q(n571)
         );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n3396), .CK(CLK), .RN(n5961), .Q(n570)
         );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n3397), .CK(CLK), .RN(RESET), .Q(n569)
         );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n3398), .CK(CLK), .RN(RESET), .Q(n568)
         );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n3399), .CK(CLK), .RN(RESET), .Q(n567)
         );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n3400), .CK(CLK), .RN(RESET), .Q(n566)
         );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n3401), .CK(CLK), .RN(RESET), .Q(n565)
         );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n3402), .CK(CLK), .RN(RESET), .Q(n564)
         );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n3403), .CK(CLK), .RN(n5954), .Q(n563)
         );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n3404), .CK(CLK), .RN(RESET), .Q(n562)
         );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n3405), .CK(CLK), .RN(n5949), .Q(n561)
         );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n3406), .CK(CLK), .RN(n5948), .Q(n560)
         );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n3407), .CK(CLK), .RN(RESET), .Q(n559)
         );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n3408), .CK(CLK), .RN(RESET), .Q(n558)
         );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n3409), .CK(CLK), .RN(RESET), .Q(n557)
         );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n3410), .CK(CLK), .RN(n5949), .Q(n556)
         );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n3411), .CK(CLK), .RN(RESET), .Q(n555)
         );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n3412), .CK(CLK), .RN(n5952), .Q(n554) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n3413), .CK(CLK), .RN(n5982), .Q(n553) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n3414), .CK(CLK), .RN(n5992), .Q(n552) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n3415), .CK(CLK), .RN(n5949), .Q(n551) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n3416), .CK(CLK), .RN(n5949), .Q(n550) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n3417), .CK(CLK), .RN(RESET), .Q(n549) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n3418), .CK(CLK), .RN(n5962), .Q(n548) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n3419), .CK(CLK), .RN(n5946), .Q(n547) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n3420), .CK(CLK), .RN(n6063), .Q(n546) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n3421), .CK(CLK), .RN(n6062), .Q(n545) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3422), .CK(CLK), .RN(RESET), .Q(n448)
         );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3423), .CK(CLK), .RN(RESET), .Q(n447)
         );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3424), .CK(CLK), .RN(n6059), .Q(n446)
         );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3425), .CK(CLK), .RN(n6062), .Q(n445)
         );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3426), .CK(CLK), .RN(n5984), .Q(n444)
         );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3427), .CK(CLK), .RN(n5983), .Q(n443)
         );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3428), .CK(CLK), .RN(RESET), .Q(n442)
         );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3429), .CK(CLK), .RN(n5946), .Q(n441)
         );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3430), .CK(CLK), .RN(n5992), .Q(n440)
         );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3431), .CK(CLK), .RN(n5958), .Q(n439)
         );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n3432), .CK(CLK), .RN(RESET), .Q(n438)
         );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n3433), .CK(CLK), .RN(n5982), .Q(n437)
         );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3434), .CK(CLK), .RN(n5983), .Q(n436)
         );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n3435), .CK(CLK), .RN(n5984), .Q(n435)
         );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3436), .CK(CLK), .RN(n5985), .Q(n434)
         );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3437), .CK(CLK), .RN(RESET), .Q(n433)
         );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3438), .CK(CLK), .RN(RESET), .Q(n432)
         );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3439), .CK(CLK), .RN(n6059), .Q(n431)
         );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3440), .CK(CLK), .RN(n6063), .Q(n430)
         );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n3441), .CK(CLK), .RN(n5993), .Q(n429)
         );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n3442), .CK(CLK), .RN(n6062), .Q(n428)
         );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3443), .CK(CLK), .RN(n6063), .Q(n427)
         );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n3444), .CK(CLK), .RN(n5992), .Q(n426) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3445), .CK(CLK), .RN(RESET), .Q(n425) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3446), .CK(CLK), .RN(RESET), .Q(n424) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3447), .CK(CLK), .RN(RESET), .Q(n423) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3448), .CK(CLK), .RN(n5954), .Q(n422) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3449), .CK(CLK), .RN(n6059), .Q(n421) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3450), .CK(CLK), .RN(RESET), .Q(n420) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3451), .CK(CLK), .RN(n5993), .Q(n419) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n3452), .CK(CLK), .RN(RESET), .Q(n418) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3453), .CK(CLK), .RN(RESET), .Q(n417) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n4157), .CK(CLK), .RN(n5946), .Q(n6236)
         );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n4156), .CK(CLK), .RN(RESET), .Q(n6237)
         );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n4155), .CK(CLK), .RN(RESET), .Q(n6238)
         );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n4154), .CK(CLK), .RN(n5955), .Q(n2270)
         );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n4153), .CK(CLK), .RN(RESET), .Q(n2265)
         );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n4152), .CK(CLK), .RN(n5962), .Q(n2260)
         );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n4151), .CK(CLK), .RN(RESET), .Q(n2255)
         );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n4150), .CK(CLK), .RN(n5992), .Q(n2250)
         );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n4149), .CK(CLK), .RN(n5983), .Q(n2245)
         );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n4148), .CK(CLK), .RN(n5954), .Q(n2240)
         );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n4147), .CK(CLK), .RN(n5955), .Q(n2235)
         );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n4146), .CK(CLK), .RN(n5956), .Q(n2230)
         );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n4145), .CK(CLK), .RN(n5957), .Q(n2225)
         );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n4144), .CK(CLK), .RN(n5958), .Q(n2220)
         );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n4143), .CK(CLK), .RN(n5959), .Q(n2215)
         );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n4142), .CK(CLK), .RN(n5960), .Q(n2210)
         );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n4141), .CK(CLK), .RN(n5961), .Q(n2205)
         );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n4140), .CK(CLK), .RN(n5962), .Q(n2200)
         );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n4139), .CK(CLK), .RN(n5963), .Q(n2195)
         );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n4138), .CK(CLK), .RN(RESET), .Q(n2190)
         );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n4137), .CK(CLK), .RN(RESET), .Q(n2185)
         );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n4136), .CK(CLK), .RN(RESET), .Q(n2180)
         );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n4135), .CK(CLK), .RN(RESET), .Q(n2175)
         );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n4134), .CK(CLK), .RN(RESET), .Q(n2170)
         );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n4133), .CK(CLK), .RN(RESET), .Q(n2165)
         );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n4132), .CK(CLK), .RN(RESET), .Q(n2160)
         );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n4131), .CK(CLK), .RN(RESET), .Q(n2155)
         );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n4130), .CK(CLK), .RN(n5974), .Q(n2150)
         );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n4129), .CK(CLK), .RN(RESET), .Q(n2145)
         );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n4128), .CK(CLK), .RN(RESET), .Q(n2140)
         );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n4127), .CK(CLK), .RN(RESET), .Q(n2135)
         );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n4126), .CK(CLK), .RN(RESET), .Q(n2130)
         );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n4125), .CK(CLK), .RN(n5946), .Q(n6239)
         );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n4124), .CK(CLK), .RN(n5985), .Q(n6240)
         );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n4123), .CK(CLK), .RN(n5984), .Q(n6241)
         );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n4122), .CK(CLK), .RN(n6063), .Q(n6242)
         );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n4121), .CK(CLK), .RN(n6062), .Q(n6243)
         );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n4120), .CK(CLK), .RN(RESET), .Q(n6244)
         );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n4119), .CK(CLK), .RN(RESET), .Q(n6245)
         );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n4118), .CK(CLK), .RN(n6059), .Q(n6246)
         );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n4117), .CK(CLK), .RN(n6063), .Q(n6247)
         );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n4116), .CK(CLK), .RN(RESET), .Q(n6248)
         );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n4115), .CK(CLK), .RN(RESET), .Q(n6249)
         );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n4114), .CK(CLK), .RN(RESET), .Q(n6250)
         );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n4113), .CK(CLK), .RN(n5974), .Q(n6251)
         );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n4112), .CK(CLK), .RN(RESET), .Q(n6252)
         );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n4111), .CK(CLK), .RN(RESET), .Q(n6253)
         );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n4110), .CK(CLK), .RN(RESET), .Q(n6254)
         );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n4109), .CK(CLK), .RN(RESET), .Q(n6255)
         );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n4108), .CK(CLK), .RN(RESET), .Q(n6256)
         );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n4107), .CK(CLK), .RN(n5982), .Q(n6257)
         );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n4106), .CK(CLK), .RN(n5983), .Q(n6258)
         );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n4105), .CK(CLK), .RN(n5984), .Q(n6259)
         );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n4104), .CK(CLK), .RN(RESET), .Q(n6260)
         );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n4103), .CK(CLK), .RN(RESET), .Q(n6261)
         );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n4102), .CK(CLK), .RN(RESET), .Q(n6262)
         );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n4101), .CK(CLK), .RN(RESET), .Q(n6263)
         );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n4100), .CK(CLK), .RN(n5974), .Q(n6264)
         );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n4099), .CK(CLK), .RN(RESET), .Q(n6265)
         );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n4098), .CK(CLK), .RN(RESET), .Q(n6266)
         );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n4097), .CK(CLK), .RN(RESET), .Q(n6267)
         );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n4096), .CK(CLK), .RN(n5955), .Q(n6268)
         );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n4095), .CK(CLK), .RN(n5948), .Q(n6269)
         );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n4094), .CK(CLK), .RN(RESET), .Q(n6270)
         );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n3454), .CK(CLK), .RN(n5982), .Q(n416)
         );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n3455), .CK(CLK), .RN(RESET), .Q(n415)
         );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n3456), .CK(CLK), .RN(n5949), .Q(n414)
         );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n3457), .CK(CLK), .RN(RESET), .Q(n413)
         );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n3458), .CK(CLK), .RN(n6059), .Q(n412)
         );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n3459), .CK(CLK), .RN(n6062), .Q(n411)
         );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n3460), .CK(CLK), .RN(n5960), .Q(n410)
         );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n3461), .CK(CLK), .RN(n5993), .Q(n409)
         );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n3462), .CK(CLK), .RN(n6063), .Q(n408)
         );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n3463), .CK(CLK), .RN(n5962), .Q(n407)
         );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n3464), .CK(CLK), .RN(n5952), .Q(n406)
         );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n3465), .CK(CLK), .RN(n6063), .Q(n405)
         );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n3466), .CK(CLK), .RN(n6062), .Q(n404)
         );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n3467), .CK(CLK), .RN(RESET), .Q(n403)
         );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n3468), .CK(CLK), .RN(RESET), .Q(n402)
         );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n3469), .CK(CLK), .RN(n6059), .Q(n401)
         );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n3470), .CK(CLK), .RN(n6062), .Q(n400)
         );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n3471), .CK(CLK), .RN(RESET), .Q(n399)
         );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n3472), .CK(CLK), .RN(n6063), .Q(n398)
         );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n3473), .CK(CLK), .RN(n6062), .Q(n397)
         );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n3474), .CK(CLK), .RN(RESET), .Q(n396)
         );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n3475), .CK(CLK), .RN(RESET), .Q(n395)
         );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n3476), .CK(CLK), .RN(RESET), .Q(n394)
         );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n3477), .CK(CLK), .RN(n5946), .Q(n393)
         );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n3478), .CK(CLK), .RN(n5963), .Q(n392)
         );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n3479), .CK(CLK), .RN(RESET), .Q(n391)
         );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n3480), .CK(CLK), .RN(n5946), .Q(n390)
         );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n3481), .CK(CLK), .RN(n5949), .Q(n389)
         );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n3482), .CK(CLK), .RN(RESET), .Q(n388)
         );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n3483), .CK(CLK), .RN(n5946), .Q(n387)
         );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n3484), .CK(CLK), .RN(RESET), .Q(n386)
         );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n3485), .CK(CLK), .RN(RESET), .Q(n385)
         );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n3486), .CK(CLK), .RN(n5946), .Q(n6271)
         );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n3487), .CK(CLK), .RN(RESET), .Q(n6272)
         );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n3488), .CK(CLK), .RN(RESET), .Q(n6273)
         );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n3489), .CK(CLK), .RN(n5974), .Q(n6274)
         );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n3490), .CK(CLK), .RN(RESET), .Q(n6275)
         );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n3491), .CK(CLK), .RN(RESET), .Q(n6276)
         );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n3492), .CK(CLK), .RN(RESET), .Q(n6277)
         );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n3493), .CK(CLK), .RN(RESET), .Q(n6278)
         );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n3494), .CK(CLK), .RN(RESET), .Q(n6279)
         );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n3495), .CK(CLK), .RN(n5982), .Q(n6280)
         );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n3496), .CK(CLK), .RN(n5983), .Q(n6281)
         );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n3497), .CK(CLK), .RN(n5984), .Q(n6282)
         );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n3498), .CK(CLK), .RN(n5985), .Q(n6283)
         );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n3499), .CK(CLK), .RN(RESET), .Q(n6284)
         );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n3500), .CK(CLK), .RN(RESET), .Q(n6285)
         );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n3501), .CK(CLK), .RN(n5959), .Q(n6286)
         );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n3502), .CK(CLK), .RN(n5992), .Q(n6287)
         );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n3503), .CK(CLK), .RN(n5952), .Q(n6288)
         );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n3504), .CK(CLK), .RN(n5954), .Q(n6289)
         );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n3505), .CK(CLK), .RN(n5955), .Q(n6290)
         );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n3506), .CK(CLK), .RN(RESET), .Q(n6291)
         );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n3507), .CK(CLK), .RN(n5960), .Q(n6292)
         );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n3508), .CK(CLK), .RN(n5992), .Q(n6293)
         );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n3509), .CK(CLK), .RN(n5956), .Q(n6294)
         );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n3510), .CK(CLK), .RN(n5957), .Q(n6295)
         );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n3511), .CK(CLK), .RN(n5958), .Q(n6296)
         );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n3512), .CK(CLK), .RN(n5959), .Q(n6297)
         );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n3513), .CK(CLK), .RN(n5960), .Q(n6298)
         );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n3514), .CK(CLK), .RN(n5961), .Q(n6299)
         );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n3515), .CK(CLK), .RN(n5962), .Q(n6300)
         );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n3516), .CK(CLK), .RN(n5963), .Q(n6301)
         );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n3517), .CK(CLK), .RN(RESET), .Q(n6302)
         );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n4093), .CK(CLK), .RN(RESET), .Q(n6303)
         );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n4092), .CK(CLK), .RN(RESET), .Q(n6304)
         );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n4091), .CK(CLK), .RN(RESET), .Q(n6305)
         );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n4090), .CK(CLK), .RN(RESET), .Q(n6306)
         );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n4089), .CK(CLK), .RN(n5974), .Q(n6307)
         );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n4088), .CK(CLK), .RN(RESET), .Q(n6308)
         );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n4087), .CK(CLK), .RN(RESET), .Q(n6309)
         );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n4086), .CK(CLK), .RN(RESET), .Q(n6310)
         );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n4085), .CK(CLK), .RN(RESET), .Q(n6311)
         );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n4084), .CK(CLK), .RN(n5952), .Q(n6312)
         );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n4083), .CK(CLK), .RN(RESET), .Q(n6313)
         );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n4082), .CK(CLK), .RN(RESET), .Q(n6314)
         );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n4081), .CK(CLK), .RN(RESET), .Q(n6315)
         );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n4080), .CK(CLK), .RN(RESET), .Q(n6316)
         );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n4079), .CK(CLK), .RN(n5946), .Q(n6317)
         );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n4078), .CK(CLK), .RN(RESET), .Q(n6318)
         );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n4077), .CK(CLK), .RN(n5946), .Q(n6319)
         );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n4076), .CK(CLK), .RN(RESET), .Q(n6320)
         );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n4075), .CK(CLK), .RN(n5946), .Q(n6321)
         );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n4074), .CK(CLK), .RN(RESET), .Q(n6322)
         );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n4073), .CK(CLK), .RN(n5946), .Q(n6323)
         );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n4072), .CK(CLK), .RN(n5949), .Q(n6324)
         );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n4071), .CK(CLK), .RN(RESET), .Q(n6325)
         );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n4070), .CK(CLK), .RN(n5946), .Q(n6326)
         );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n4069), .CK(CLK), .RN(RESET), .Q(n6327)
         );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n4068), .CK(CLK), .RN(RESET), .Q(n6328)
         );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n4067), .CK(CLK), .RN(RESET), .Q(n6329)
         );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n4066), .CK(CLK), .RN(RESET), .Q(n6330)
         );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n4065), .CK(CLK), .RN(RESET), .Q(n6331)
         );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n4064), .CK(CLK), .RN(RESET), .Q(n6332)
         );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n4063), .CK(CLK), .RN(RESET), .Q(n6333)
         );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n4062), .CK(CLK), .RN(RESET), .Q(n6334)
         );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n4061), .CK(CLK), .RN(RESET), .Q(n2382)
         );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n4060), .CK(CLK), .RN(n5974), .Q(n2379)
         );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n4059), .CK(CLK), .RN(RESET), .Q(n2376)
         );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n4058), .CK(CLK), .RN(RESET), .Q(n2373)
         );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n4057), .CK(CLK), .RN(RESET), .Q(n2370)
         );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n4056), .CK(CLK), .RN(RESET), .Q(n2367)
         );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n4055), .CK(CLK), .RN(RESET), .Q(n2364)
         );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n4054), .CK(CLK), .RN(RESET), .Q(n2361)
         );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n4053), .CK(CLK), .RN(RESET), .Q(n2358)
         );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n4052), .CK(CLK), .RN(RESET), .Q(n2355)
         );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n4051), .CK(CLK), .RN(RESET), .Q(n2352)
         );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n4050), .CK(CLK), .RN(n5974), .Q(n6335)
         );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n4049), .CK(CLK), .RN(RESET), .Q(n6336)
         );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n4048), .CK(CLK), .RN(RESET), .Q(n6337)
         );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n4047), .CK(CLK), .RN(n5983), .Q(n6338)
         );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n4046), .CK(CLK), .RN(n5984), .Q(n6339)
         );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n4045), .CK(CLK), .RN(n5985), .Q(n6340)
         );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n4044), .CK(CLK), .RN(RESET), .Q(n6341)
         );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n4043), .CK(CLK), .RN(RESET), .Q(n6342)
         );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n4042), .CK(CLK), .RN(RESET), .Q(n6343)
         );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n4041), .CK(CLK), .RN(n5982), .Q(n6344)
         );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n4040), .CK(CLK), .RN(n5983), .Q(n6345)
         );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n4039), .CK(CLK), .RN(n5984), .Q(n6346)
         );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n4038), .CK(CLK), .RN(n5985), .Q(n6347)
         );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n4037), .CK(CLK), .RN(RESET), .Q(n6348)
         );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n4036), .CK(CLK), .RN(RESET), .Q(n6349)
         );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n4035), .CK(CLK), .RN(RESET), .Q(n6350)
         );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n4034), .CK(CLK), .RN(n5974), .Q(n6351)
         );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n4033), .CK(CLK), .RN(RESET), .Q(n6352)
         );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n4032), .CK(CLK), .RN(RESET), .Q(n6353)
         );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n4031), .CK(CLK), .RN(RESET), .Q(n6354)
         );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n4030), .CK(CLK), .RN(RESET), .Q(n6355)
         );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n3518), .CK(CLK), .RN(n5961), .Q(n704)
         );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n3519), .CK(CLK), .RN(n5992), .Q(n703)
         );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n3520), .CK(CLK), .RN(RESET), .Q(n702)
         );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n3521), .CK(CLK), .RN(RESET), .Q(n701)
         );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n3522), .CK(CLK), .RN(n5952), .Q(n700)
         );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n3523), .CK(CLK), .RN(n5954), .Q(n699)
         );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n3524), .CK(CLK), .RN(n5955), .Q(n698)
         );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n3525), .CK(CLK), .RN(n5956), .Q(n697)
         );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n3526), .CK(CLK), .RN(n6062), .Q(n696)
         );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n3527), .CK(CLK), .RN(n5993), .Q(n695)
         );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n3528), .CK(CLK), .RN(n5952), .Q(n694)
         );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n3529), .CK(CLK), .RN(n6059), .Q(n693)
         );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n3530), .CK(CLK), .RN(RESET), .Q(n692)
         );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n3531), .CK(CLK), .RN(n5956), .Q(n691)
         );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n3532), .CK(CLK), .RN(RESET), .Q(n690)
         );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n3533), .CK(CLK), .RN(n5957), .Q(n689)
         );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n3534), .CK(CLK), .RN(n5958), .Q(n688)
         );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n3535), .CK(CLK), .RN(n5959), .Q(n687)
         );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n3536), .CK(CLK), .RN(n5960), .Q(n686)
         );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n3537), .CK(CLK), .RN(n5961), .Q(n685)
         );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n3538), .CK(CLK), .RN(n5962), .Q(n684)
         );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n3539), .CK(CLK), .RN(n5963), .Q(n683)
         );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n3540), .CK(CLK), .RN(RESET), .Q(n682)
         );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n3541), .CK(CLK), .RN(RESET), .Q(n681)
         );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n3542), .CK(CLK), .RN(RESET), .Q(n680)
         );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n3543), .CK(CLK), .RN(RESET), .Q(n679)
         );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n3544), .CK(CLK), .RN(RESET), .Q(n678)
         );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n3545), .CK(CLK), .RN(n6059), .Q(n677)
         );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n3546), .CK(CLK), .RN(n5948), .Q(n676)
         );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n3547), .CK(CLK), .RN(RESET), .Q(n675)
         );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n3548), .CK(CLK), .RN(RESET), .Q(n674)
         );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n3549), .CK(CLK), .RN(n6059), .Q(n673)
         );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n3550), .CK(CLK), .RN(n5948), .Q(n6356)
         );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n3551), .CK(CLK), .RN(RESET), .Q(n6357)
         );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n3552), .CK(CLK), .RN(RESET), .Q(n6358)
         );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n3553), .CK(CLK), .RN(n6059), .Q(n6359)
         );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n3554), .CK(CLK), .RN(n5948), .Q(n6360)
         );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n3555), .CK(CLK), .RN(RESET), .Q(n6361)
         );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n3556), .CK(CLK), .RN(n5946), .Q(n6362)
         );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n3557), .CK(CLK), .RN(n5957), .Q(n6363)
         );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n3558), .CK(CLK), .RN(n5958), .Q(n6364)
         );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n3559), .CK(CLK), .RN(n5959), .Q(n6365)
         );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n3560), .CK(CLK), .RN(n5960), .Q(n6366)
         );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n3561), .CK(CLK), .RN(n5961), .Q(n6367)
         );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n3562), .CK(CLK), .RN(n5962), .Q(n6368)
         );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n3563), .CK(CLK), .RN(n5963), .Q(n6369)
         );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n3564), .CK(CLK), .RN(RESET), .Q(n6370)
         );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n3565), .CK(CLK), .RN(n5993), .Q(n6371)
         );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n3566), .CK(CLK), .RN(n5958), .Q(n6372)
         );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n3567), .CK(CLK), .RN(n5959), .Q(n6373)
         );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n3568), .CK(CLK), .RN(n5960), .Q(n6374)
         );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n3569), .CK(CLK), .RN(n5961), .Q(n6375)
         );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n3570), .CK(CLK), .RN(n5962), .Q(n6376)
         );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n3571), .CK(CLK), .RN(n5963), .Q(n6377)
         );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n3572), .CK(CLK), .RN(RESET), .Q(n6378)
         );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n3573), .CK(CLK), .RN(n5993), .Q(n6379)
         );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n3574), .CK(CLK), .RN(n5963), .Q(n6380)
         );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n3575), .CK(CLK), .RN(n5993), .Q(n6381)
         );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n3576), .CK(CLK), .RN(n5954), .Q(n6382)
         );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n3577), .CK(CLK), .RN(n5952), .Q(n6383)
         );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n3578), .CK(CLK), .RN(RESET), .Q(n6384)
         );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n3579), .CK(CLK), .RN(RESET), .Q(n6385)
         );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n3580), .CK(CLK), .RN(RESET), .Q(n6386)
         );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n3581), .CK(CLK), .RN(RESET), .Q(n6387)
         );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n4029), .CK(CLK), .RN(RESET), .Q(n6388)
         );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n4028), .CK(CLK), .RN(RESET), .Q(n6389)
         );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n4027), .CK(CLK), .RN(RESET), .Q(n6390)
         );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n4026), .CK(CLK), .RN(RESET), .Q(n6391)
         );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n4025), .CK(CLK), .RN(RESET), .Q(n6392)
         );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n4024), .CK(CLK), .RN(RESET), .Q(n6393)
         );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n4023), .CK(CLK), .RN(RESET), .Q(n6394)
         );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n4022), .CK(CLK), .RN(RESET), .Q(n6395)
         );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n4021), .CK(CLK), .RN(RESET), .Q(n6396)
         );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n4020), .CK(CLK), .RN(RESET), .Q(n6397)
         );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n4019), .CK(CLK), .RN(RESET), .Q(n6398)
         );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n4018), .CK(CLK), .RN(RESET), .Q(n6399)
         );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n4017), .CK(CLK), .RN(RESET), .Q(n6400)
         );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n4016), .CK(CLK), .RN(RESET), .Q(n6401)
         );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n4015), .CK(CLK), .RN(RESET), .Q(n6402)
         );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n4014), .CK(CLK), .RN(RESET), .Q(n6403)
         );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n4013), .CK(CLK), .RN(RESET), .Q(n6404)
         );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n4012), .CK(CLK), .RN(RESET), .Q(n6405)
         );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n4011), .CK(CLK), .RN(RESET), .Q(n6406)
         );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n4010), .CK(CLK), .RN(RESET), .Q(n6407)
         );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n4009), .CK(CLK), .RN(n5963), .Q(n6408)
         );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n4008), .CK(CLK), .RN(n5992), .Q(n6409)
         );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n4007), .CK(CLK), .RN(n5952), .Q(n6410)
         );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n4006), .CK(CLK), .RN(RESET), .Q(n6411)
         );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n4005), .CK(CLK), .RN(RESET), .Q(n6412)
         );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n4004), .CK(CLK), .RN(RESET), .Q(n6413)
         );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n4003), .CK(CLK), .RN(RESET), .Q(n6414)
         );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n4002), .CK(CLK), .RN(RESET), .Q(n6415)
         );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n4001), .CK(CLK), .RN(n5954), .Q(n6416)
         );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n4000), .CK(CLK), .RN(n5955), .Q(n6417)
         );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3999), .CK(CLK), .RN(n5956), .Q(n6418)
         );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3998), .CK(CLK), .RN(RESET), .Q(n6419)
         );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3790), .CK(CLK), .RN(n5957), .Q(n6420)
         );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3789), .CK(CLK), .RN(n5958), .Q(n6421)
         );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3788), .CK(CLK), .RN(n5959), .Q(n6422)
         );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3787), .CK(CLK), .RN(n5960), .Q(n6423)
         );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3786), .CK(CLK), .RN(n5961), .Q(n6424)
         );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3785), .CK(CLK), .RN(n5962), .Q(n6425)
         );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3784), .CK(CLK), .RN(n5963), .Q(n6426)
         );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3783), .CK(CLK), .RN(RESET), .Q(n6427)
         );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3782), .CK(CLK), .RN(n6059), .Q(n6428)
         );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3781), .CK(CLK), .RN(n5948), .Q(n6429)
         );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3780), .CK(CLK), .RN(n6063), .Q(n6430)
         );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3779), .CK(CLK), .RN(n6062), .Q(n6431)
         );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3778), .CK(CLK), .RN(RESET), .Q(n6432)
         );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3777), .CK(CLK), .RN(RESET), .Q(n6433)
         );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3776), .CK(CLK), .RN(n6059), .Q(n6434)
         );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3775), .CK(CLK), .RN(n5948), .Q(n6435)
         );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3774), .CK(CLK), .RN(n6063), .Q(n6436)
         );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3165), .CK(CLK), .RN(n6062), .Q(n6437)
         );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3164), .CK(CLK), .RN(n5993), .Q(n6438)
         );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3163), .CK(CLK), .RN(n5993), .Q(n6439)
         );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3162), .CK(CLK), .RN(n5993), .Q(n6440)
         );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3161), .CK(CLK), .RN(n5993), .Q(n6441)
         );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3160), .CK(CLK), .RN(n5993), .Q(n6442)
         );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3159), .CK(CLK), .RN(n5993), .Q(n6443)
         );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3158), .CK(CLK), .RN(n5993), .Q(n6444)
         );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3157), .CK(CLK), .RN(n5993), .Q(n6445)
         );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3156), .CK(CLK), .RN(n5993), .Q(n6446)
         );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3155), .CK(CLK), .RN(n5993), .Q(n6447)
         );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3154), .CK(CLK), .RN(n5993), .Q(n6448)
         );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3153), .CK(CLK), .RN(n5992), .Q(n6449)
         );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3152), .CK(CLK), .RN(n5992), .Q(n6450)
         );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3151), .CK(CLK), .RN(n5992), .Q(n6451)
         );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n3582), .CK(CLK), .RN(n5992), .Q(n736)
         );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n3583), .CK(CLK), .RN(n5992), .Q(n735)
         );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n3584), .CK(CLK), .RN(n5992), .Q(n734)
         );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n3585), .CK(CLK), .RN(n5992), .Q(n733)
         );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n3586), .CK(CLK), .RN(n5992), .Q(n732)
         );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n3587), .CK(CLK), .RN(n5992), .Q(n731)
         );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n3588), .CK(CLK), .RN(n5992), .Q(n730)
         );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n3589), .CK(CLK), .RN(n5992), .Q(n729)
         );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n3590), .CK(CLK), .RN(n5955), .Q(n728)
         );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n3591), .CK(CLK), .RN(n5956), .Q(n727)
         );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n3592), .CK(CLK), .RN(n5957), .Q(n726)
         );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n3593), .CK(CLK), .RN(n5958), .Q(n725)
         );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n3594), .CK(CLK), .RN(n5959), .Q(n724)
         );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n3595), .CK(CLK), .RN(n5960), .Q(n723)
         );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n3596), .CK(CLK), .RN(n5961), .Q(n722)
         );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n3597), .CK(CLK), .RN(n5962), .Q(n721)
         );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n3598), .CK(CLK), .RN(n5963), .Q(n720)
         );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n3599), .CK(CLK), .RN(n5954), .Q(n719)
         );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n3600), .CK(CLK), .RN(n5955), .Q(n718)
         );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n3601), .CK(CLK), .RN(n5948), .Q(n717)
         );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n3602), .CK(CLK), .RN(n5948), .Q(n716)
         );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n3603), .CK(CLK), .RN(n6063), .Q(n715)
         );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n3604), .CK(CLK), .RN(n5948), .Q(n714)
         );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n3605), .CK(CLK), .RN(RESET), .Q(n713)
         );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n3606), .CK(CLK), .RN(n5948), .Q(n712)
         );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n3607), .CK(CLK), .RN(n5946), .Q(n711)
         );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n3608), .CK(CLK), .RN(n5946), .Q(n710)
         );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n3609), .CK(CLK), .RN(n5948), .Q(n709)
         );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n3610), .CK(CLK), .RN(n6063), .Q(n708)
         );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n3611), .CK(CLK), .RN(n6062), .Q(n707)
         );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n3612), .CK(CLK), .RN(RESET), .Q(n706)
         );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n3613), .CK(CLK), .RN(RESET), .Q(n705)
         );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n3614), .CK(CLK), .RN(RESET), .Q(n544)
         );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n3615), .CK(CLK), .RN(RESET), .Q(n543)
         );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n3616), .CK(CLK), .RN(n6059), .Q(n542)
         );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n3617), .CK(CLK), .RN(RESET), .Q(n541)
         );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n3618), .CK(CLK), .RN(RESET), .Q(n540)
         );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n3619), .CK(CLK), .RN(n6059), .Q(n539)
         );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n3620), .CK(CLK), .RN(RESET), .Q(n538)
         );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n3621), .CK(CLK), .RN(n6059), .Q(n537)
         );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n3622), .CK(CLK), .RN(RESET), .Q(n536)
         );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n3623), .CK(CLK), .RN(n5948), .Q(n535)
         );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n3624), .CK(CLK), .RN(n5946), .Q(n534)
         );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n3625), .CK(CLK), .RN(n5948), .Q(n533)
         );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n3626), .CK(CLK), .RN(n5948), .Q(n532)
         );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n3627), .CK(CLK), .RN(RESET), .Q(n531)
         );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n3628), .CK(CLK), .RN(RESET), .Q(n530)
         );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n3629), .CK(CLK), .RN(n6063), .Q(n529)
         );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n3630), .CK(CLK), .RN(n5948), .Q(n528)
         );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n3631), .CK(CLK), .RN(RESET), .Q(n527)
         );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n3632), .CK(CLK), .RN(RESET), .Q(n526)
         );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n3633), .CK(CLK), .RN(n5948), .Q(n525)
         );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n3634), .CK(CLK), .RN(RESET), .Q(n524)
         );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n3635), .CK(CLK), .RN(RESET), .Q(n523)
         );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n3636), .CK(CLK), .RN(RESET), .Q(n522)
         );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n3637), .CK(CLK), .RN(RESET), .Q(n521)
         );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n3638), .CK(CLK), .RN(RESET), .Q(n520)
         );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n3639), .CK(CLK), .RN(RESET), .Q(n519)
         );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n3640), .CK(CLK), .RN(RESET), .Q(n518)
         );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n3641), .CK(CLK), .RN(RESET), .Q(n517)
         );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n3642), .CK(CLK), .RN(RESET), .Q(n516)
         );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n3643), .CK(CLK), .RN(RESET), .Q(n515)
         );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n3644), .CK(CLK), .RN(RESET), .Q(n514)
         );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n3645), .CK(CLK), .RN(RESET), .Q(n513)
         );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3886), .CK(CLK), .RN(RESET), .Q(n6452)
         );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3885), .CK(CLK), .RN(RESET), .Q(n6453)
         );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3884), .CK(CLK), .RN(RESET), .Q(n6454)
         );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3883), .CK(CLK), .RN(RESET), .Q(n6455)
         );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3882), .CK(CLK), .RN(RESET), .Q(n6456)
         );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3881), .CK(CLK), .RN(RESET), .Q(n6457)
         );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3880), .CK(CLK), .RN(RESET), .Q(n6458)
         );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3879), .CK(CLK), .RN(RESET), .Q(n6459)
         );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3878), .CK(CLK), .RN(RESET), .Q(n6460)
         );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3877), .CK(CLK), .RN(RESET), .Q(n6461)
         );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3876), .CK(CLK), .RN(n5985), .Q(n6462)
         );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3875), .CK(CLK), .RN(n5985), .Q(n6463)
         );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3874), .CK(CLK), .RN(n5985), .Q(n6464)
         );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3873), .CK(CLK), .RN(n5985), .Q(n6465)
         );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3872), .CK(CLK), .RN(n5985), .Q(n6466)
         );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3871), .CK(CLK), .RN(n5985), .Q(n6467)
         );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3870), .CK(CLK), .RN(n5985), .Q(n6468)
         );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3805), .CK(CLK), .RN(n5985), .Q(n6469)
         );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3804), .CK(CLK), .RN(n5985), .Q(n6470)
         );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3803), .CK(CLK), .RN(n5985), .Q(n6471)
         );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3802), .CK(CLK), .RN(n5985), .Q(n6472)
         );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3801), .CK(CLK), .RN(n5984), .Q(n6473)
         );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3800), .CK(CLK), .RN(n5984), .Q(n6474)
         );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3799), .CK(CLK), .RN(n5984), .Q(n6475)
         );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3798), .CK(CLK), .RN(n5984), .Q(n6476)
         );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3797), .CK(CLK), .RN(n5984), .Q(n6477)
         );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3796), .CK(CLK), .RN(n5984), .Q(n6478)
         );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3795), .CK(CLK), .RN(n5984), .Q(n6479)
         );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3794), .CK(CLK), .RN(n5984), .Q(n6480)
         );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3793), .CK(CLK), .RN(n5984), .Q(n6481)
         );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3792), .CK(CLK), .RN(n5984), .Q(n6482)
         );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3791), .CK(CLK), .RN(n5984), .Q(n6483)
         );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3918), .CK(CLK), .RN(n5983), .Q(n6484), 
        .QN(n1423) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3917), .CK(CLK), .RN(n5983), .Q(n6485), 
        .QN(n1424) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n3916), .CK(CLK), .RN(n5983), .Q(n6486), 
        .QN(n1425) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n3915), .CK(CLK), .RN(n5983), .Q(n6487), 
        .QN(n1426) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3914), .CK(CLK), .RN(n5983), .Q(n6488), 
        .QN(n1427) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3913), .CK(CLK), .RN(n5983), .Q(n6489), 
        .QN(n1428) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3912), .CK(CLK), .RN(n5983), .Q(n6490), 
        .QN(n1429) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n3911), .CK(CLK), .RN(n5983), .Q(n6491), 
        .QN(n1430) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3910), .CK(CLK), .RN(n5983), .Q(n6492), 
        .QN(n1431) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n3909), .CK(CLK), .RN(n5983), .Q(n6493), 
        .QN(n1432) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n3908), .CK(CLK), .RN(n5983), .Q(n6494), 
        .QN(n1433) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n3907), .CK(CLK), .RN(n5982), .Q(n6495), 
        .QN(n1434) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3906), .CK(CLK), .RN(n5982), .Q(n6496), 
        .QN(n1435) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n3905), .CK(CLK), .RN(n5982), .Q(n6497), 
        .QN(n1436) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3904), .CK(CLK), .RN(n5982), .Q(n6498), 
        .QN(n1437) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3903), .CK(CLK), .RN(n5982), .Q(n6499), 
        .QN(n1438) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3902), .CK(CLK), .RN(n5982), .Q(n6500), 
        .QN(n1439) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3901), .CK(CLK), .RN(n5982), .Q(n6501), 
        .QN(n1440) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3900), .CK(CLK), .RN(n5982), .Q(n6502), 
        .QN(n1441) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n3899), .CK(CLK), .RN(n5982), .Q(n6503), 
        .QN(n1442) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n3898), .CK(CLK), .RN(n5982), .Q(n6504), 
        .QN(n1443) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3897), .CK(CLK), .RN(n5982), .Q(n6505), 
        .QN(n1444) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3896), .CK(CLK), .RN(RESET), .Q(n6506), 
        .QN(n1445) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3895), .CK(CLK), .RN(RESET), .Q(n6507), 
        .QN(n1446) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3894), .CK(CLK), .RN(RESET), .Q(n6508), 
        .QN(n1447) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3893), .CK(CLK), .RN(RESET), .Q(n6509), 
        .QN(n1448) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n3892), .CK(CLK), .RN(RESET), .Q(n6510), 
        .QN(n1449) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3891), .CK(CLK), .RN(RESET), .Q(n6511), 
        .QN(n1450) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3890), .CK(CLK), .RN(RESET), .Q(n6512), 
        .QN(n1451) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3889), .CK(CLK), .RN(RESET), .Q(n6513), 
        .QN(n1452) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3888), .CK(CLK), .RN(RESET), .Q(n6514), 
        .QN(n1453) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3887), .CK(CLK), .RN(RESET), .Q(n6515), 
        .QN(n1454) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3118), .CK(CLK), .RN(RESET), .Q(n6516)
         );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n3117), .CK(CLK), .RN(RESET), .Q(n6517)
         );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n3116), .CK(CLK), .RN(RESET), .Q(n6518)
         );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n3115), .CK(CLK), .RN(RESET), .Q(n6519)
         );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n3114), .CK(CLK), .RN(RESET), .Q(n6520)
         );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n3113), .CK(CLK), .RN(RESET), .Q(n6521)
         );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n3112), .CK(CLK), .RN(RESET), .Q(n6522)
         );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n3111), .CK(CLK), .RN(RESET), .Q(n6523)
         );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n3110), .CK(CLK), .RN(RESET), .Q(n6524)
         );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n3109), .CK(CLK), .RN(RESET), .Q(n6525)
         );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n3108), .CK(CLK), .RN(RESET), .Q(n6526)
         );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n3107), .CK(CLK), .RN(RESET), .Q(n6527)
         );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n3106), .CK(CLK), .RN(RESET), .Q(n6528)
         );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n3105), .CK(CLK), .RN(RESET), .Q(n6529)
         );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n3104), .CK(CLK), .RN(RESET), .Q(n6530)
         );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n3103), .CK(CLK), .RN(RESET), .Q(n6531)
         );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n3102), .CK(CLK), .RN(RESET), .Q(n6532)
         );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n3101), .CK(CLK), .RN(RESET), .Q(n6533)
         );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n3100), .CK(CLK), .RN(RESET), .Q(n6534)
         );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n3099), .CK(CLK), .RN(RESET), .Q(n6535)
         );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n3098), .CK(CLK), .RN(RESET), .Q(n6536)
         );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n3097), .CK(CLK), .RN(RESET), .Q(n6537)
         );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n3096), .CK(CLK), .RN(RESET), .Q(n6538)
         );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n3095), .CK(CLK), .RN(RESET), .Q(n6539)
         );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n3094), .CK(CLK), .RN(RESET), .Q(n6540)
         );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n3093), .CK(CLK), .RN(RESET), .Q(n6541)
         );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n3092), .CK(CLK), .RN(RESET), .Q(n6542)
         );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n3091), .CK(CLK), .RN(RESET), .Q(n6543)
         );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3090), .CK(CLK), .RN(RESET), .Q(n6544)
         );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3089), .CK(CLK), .RN(RESET), .Q(n6545)
         );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3088), .CK(CLK), .RN(RESET), .Q(n6546)
         );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3087), .CK(CLK), .RN(RESET), .Q(n6547)
         );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3869), .CK(CLK), .RN(RESET), .Q(n2830)
         );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3868), .CK(CLK), .RN(RESET), .Q(n2829)
         );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3867), .CK(CLK), .RN(RESET), .Q(n2828)
         );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3866), .CK(CLK), .RN(RESET), .Q(n2827)
         );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3865), .CK(CLK), .RN(RESET), .Q(n2826)
         );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3864), .CK(CLK), .RN(RESET), .Q(n2825)
         );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3863), .CK(CLK), .RN(RESET), .Q(n2824)
         );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3862), .CK(CLK), .RN(RESET), .Q(n2823)
         );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3861), .CK(CLK), .RN(RESET), .Q(n2822)
         );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3860), .CK(CLK), .RN(RESET), .Q(n2821)
         );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3859), .CK(CLK), .RN(RESET), .Q(n2820)
         );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3858), .CK(CLK), .RN(RESET), .Q(n2819)
         );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3857), .CK(CLK), .RN(RESET), .Q(n2818)
         );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3856), .CK(CLK), .RN(RESET), .Q(n2817)
         );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3855), .CK(CLK), .RN(RESET), .Q(n2816)
         );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3854), .CK(CLK), .RN(RESET), .Q(n2815)
         );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3853), .CK(CLK), .RN(RESET), .Q(n2814)
         );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3852), .CK(CLK), .RN(RESET), .Q(n2813)
         );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3851), .CK(CLK), .RN(RESET), .Q(n2812)
         );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3850), .CK(CLK), .RN(RESET), .Q(n2811)
         );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3849), .CK(CLK), .RN(RESET), .Q(n2810)
         );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3848), .CK(CLK), .RN(RESET), .Q(n2809)
         );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3847), .CK(CLK), .RN(RESET), .Q(n2808)
         );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3846), .CK(CLK), .RN(RESET), .Q(n2807)
         );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3845), .CK(CLK), .RN(RESET), .Q(n6548)
         );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3844), .CK(CLK), .RN(RESET), .Q(n6549)
         );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3843), .CK(CLK), .RN(RESET), .Q(n6550)
         );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3842), .CK(CLK), .RN(RESET), .Q(n6551)
         );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3841), .CK(CLK), .RN(RESET), .Q(n6552)
         );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3840), .CK(CLK), .RN(RESET), .Q(n6553)
         );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3839), .CK(CLK), .RN(RESET), .Q(n6554)
         );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3838), .CK(CLK), .RN(RESET), .Q(n6555)
         );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n3646), .CK(CLK), .RN(RESET), .Q(n512)
         );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n3647), .CK(CLK), .RN(RESET), .Q(n511)
         );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n3648), .CK(CLK), .RN(RESET), .Q(n510)
         );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n3649), .CK(CLK), .RN(n5974), .Q(n509)
         );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n3650), .CK(CLK), .RN(n5974), .Q(n508)
         );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n3651), .CK(CLK), .RN(n5974), .Q(n507)
         );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n3652), .CK(CLK), .RN(n5974), .Q(n506)
         );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n3653), .CK(CLK), .RN(n5974), .Q(n505)
         );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n3654), .CK(CLK), .RN(n5974), .Q(n504)
         );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n3655), .CK(CLK), .RN(n5974), .Q(n503)
         );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n3656), .CK(CLK), .RN(n5974), .Q(n502)
         );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n3657), .CK(CLK), .RN(n5974), .Q(n501)
         );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n3658), .CK(CLK), .RN(n5974), .Q(n500)
         );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n3659), .CK(CLK), .RN(n5974), .Q(n499)
         );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n3660), .CK(CLK), .RN(RESET), .Q(n498)
         );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n3661), .CK(CLK), .RN(RESET), .Q(n497)
         );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n3662), .CK(CLK), .RN(RESET), .Q(n496)
         );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n3663), .CK(CLK), .RN(RESET), .Q(n495)
         );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n3664), .CK(CLK), .RN(RESET), .Q(n494)
         );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n3665), .CK(CLK), .RN(RESET), .Q(n493)
         );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n3666), .CK(CLK), .RN(RESET), .Q(n492)
         );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n3667), .CK(CLK), .RN(RESET), .Q(n491)
         );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n3668), .CK(CLK), .RN(RESET), .Q(n490)
         );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n3669), .CK(CLK), .RN(RESET), .Q(n489)
         );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n3670), .CK(CLK), .RN(RESET), .Q(n488)
         );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n3671), .CK(CLK), .RN(RESET), .Q(n487)
         );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n3672), .CK(CLK), .RN(RESET), .Q(n486)
         );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n3673), .CK(CLK), .RN(RESET), .Q(n485)
         );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n3674), .CK(CLK), .RN(RESET), .Q(n484)
         );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n3675), .CK(CLK), .RN(RESET), .Q(n483)
         );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n3676), .CK(CLK), .RN(RESET), .Q(n482)
         );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n3677), .CK(CLK), .RN(RESET), .Q(n481)
         );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n3678), .CK(CLK), .RN(RESET), .Q(n672)
         );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n3679), .CK(CLK), .RN(RESET), .Q(n671)
         );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n3680), .CK(CLK), .RN(RESET), .Q(n670)
         );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n3681), .CK(CLK), .RN(RESET), .Q(n669)
         );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n3682), .CK(CLK), .RN(RESET), .Q(n668)
         );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n3683), .CK(CLK), .RN(RESET), .Q(n667)
         );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n3684), .CK(CLK), .RN(RESET), .Q(n666)
         );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n3685), .CK(CLK), .RN(RESET), .Q(n665)
         );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n3686), .CK(CLK), .RN(RESET), .Q(n664)
         );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n3687), .CK(CLK), .RN(RESET), .Q(n663)
         );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n3688), .CK(CLK), .RN(RESET), .Q(n662)
         );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n3689), .CK(CLK), .RN(RESET), .Q(n661)
         );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n3690), .CK(CLK), .RN(RESET), .Q(n660)
         );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n3691), .CK(CLK), .RN(RESET), .Q(n659)
         );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n3692), .CK(CLK), .RN(RESET), .Q(n658)
         );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n3693), .CK(CLK), .RN(RESET), .Q(n657)
         );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n3694), .CK(CLK), .RN(RESET), .Q(n656)
         );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n3695), .CK(CLK), .RN(RESET), .Q(n655)
         );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n3696), .CK(CLK), .RN(RESET), .Q(n654)
         );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n3697), .CK(CLK), .RN(RESET), .Q(n653)
         );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n3698), .CK(CLK), .RN(RESET), .Q(n652)
         );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n3699), .CK(CLK), .RN(RESET), .Q(n651)
         );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n3700), .CK(CLK), .RN(RESET), .Q(n650)
         );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n3701), .CK(CLK), .RN(RESET), .Q(n649)
         );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n3702), .CK(CLK), .RN(RESET), .Q(n648)
         );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n3703), .CK(CLK), .RN(RESET), .Q(n647)
         );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n3704), .CK(CLK), .RN(RESET), .Q(n646)
         );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n3705), .CK(CLK), .RN(RESET), .Q(n645)
         );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n3706), .CK(CLK), .RN(RESET), .Q(n644)
         );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n3707), .CK(CLK), .RN(RESET), .Q(n643)
         );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n3708), .CK(CLK), .RN(RESET), .Q(n642)
         );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n3709), .CK(CLK), .RN(RESET), .Q(n641)
         );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3837), .CK(CLK), .RN(RESET), .Q(n6556)
         );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3836), .CK(CLK), .RN(RESET), .Q(n6557)
         );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3835), .CK(CLK), .RN(RESET), .Q(n6558)
         );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3834), .CK(CLK), .RN(RESET), .Q(n6559)
         );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3833), .CK(CLK), .RN(RESET), .Q(n6560)
         );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3832), .CK(CLK), .RN(RESET), .Q(n6561)
         );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3831), .CK(CLK), .RN(RESET), .Q(n6562)
         );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3830), .CK(CLK), .RN(RESET), .Q(n6563)
         );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3829), .CK(CLK), .RN(RESET), .Q(n6564)
         );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3828), .CK(CLK), .RN(RESET), .Q(n6565)
         );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3827), .CK(CLK), .RN(RESET), .Q(n6566)
         );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3826), .CK(CLK), .RN(RESET), .Q(n6567)
         );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3825), .CK(CLK), .RN(RESET), .Q(n6568)
         );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3824), .CK(CLK), .RN(RESET), .Q(n6569)
         );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3823), .CK(CLK), .RN(RESET), .Q(n6570)
         );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3822), .CK(CLK), .RN(RESET), .Q(n6571)
         );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3821), .CK(CLK), .RN(RESET), .Q(n6572)
         );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3820), .CK(CLK), .RN(RESET), .Q(n6573)
         );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3819), .CK(CLK), .RN(RESET), .Q(n6574)
         );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3818), .CK(CLK), .RN(RESET), .Q(n6575)
         );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3817), .CK(CLK), .RN(RESET), .Q(n6576)
         );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3816), .CK(CLK), .RN(RESET), .Q(n6577)
         );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3815), .CK(CLK), .RN(RESET), .Q(n6578)
         );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3814), .CK(CLK), .RN(RESET), .Q(n6579)
         );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3813), .CK(CLK), .RN(RESET), .Q(n6580)
         );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3812), .CK(CLK), .RN(RESET), .Q(n6581)
         );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3811), .CK(CLK), .RN(RESET), .Q(n6582)
         );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3810), .CK(CLK), .RN(RESET), .Q(n6583)
         );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3809), .CK(CLK), .RN(RESET), .Q(n6584)
         );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3808), .CK(CLK), .RN(RESET), .Q(n6585)
         );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3807), .CK(CLK), .RN(RESET), .Q(n6586)
         );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3806), .CK(CLK), .RN(RESET), .Q(n6587)
         );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3150), .CK(CLK), .RN(RESET), .Q(n6588)
         );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3149), .CK(CLK), .RN(RESET), .Q(n6589)
         );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3148), .CK(CLK), .RN(RESET), .Q(n6590)
         );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3147), .CK(CLK), .RN(RESET), .Q(n6591)
         );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3146), .CK(CLK), .RN(RESET), .Q(n6592)
         );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3145), .CK(CLK), .RN(RESET), .Q(n6593)
         );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3144), .CK(CLK), .RN(RESET), .Q(n6594)
         );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3143), .CK(CLK), .RN(RESET), .Q(n6595)
         );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3142), .CK(CLK), .RN(RESET), .Q(n6596)
         );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3141), .CK(CLK), .RN(RESET), .Q(n6597)
         );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3140), .CK(CLK), .RN(RESET), .Q(n6598)
         );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3139), .CK(CLK), .RN(RESET), .Q(n6599)
         );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3138), .CK(CLK), .RN(RESET), .Q(n6600)
         );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3137), .CK(CLK), .RN(RESET), .Q(n6601)
         );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3136), .CK(CLK), .RN(RESET), .Q(n6602)
         );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3135), .CK(CLK), .RN(RESET), .Q(n6603)
         );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3134), .CK(CLK), .RN(RESET), .Q(n6604)
         );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3133), .CK(CLK), .RN(RESET), .Q(n6605)
         );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3132), .CK(CLK), .RN(RESET), .Q(n6606)
         );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3131), .CK(CLK), .RN(RESET), .Q(n6607)
         );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3130), .CK(CLK), .RN(RESET), .Q(n6608)
         );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3129), .CK(CLK), .RN(RESET), .Q(n6609)
         );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3128), .CK(CLK), .RN(RESET), .Q(n6610)
         );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3127), .CK(CLK), .RN(RESET), .Q(n6611)
         );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3126), .CK(CLK), .RN(RESET), .Q(n6612)
         );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3125), .CK(CLK), .RN(RESET), .Q(n6613)
         );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3124), .CK(CLK), .RN(RESET), .Q(n6614)
         );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3123), .CK(CLK), .RN(RESET), .Q(n6615)
         );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3122), .CK(CLK), .RN(n5963), .Q(n6616)
         );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3121), .CK(CLK), .RN(n5963), .Q(n6617)
         );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3120), .CK(CLK), .RN(n5963), .Q(n6618)
         );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3119), .CK(CLK), .RN(n5963), .Q(n6619)
         );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n3710), .CK(CLK), .RN(n5963), .Q(n384)
         );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n3711), .CK(CLK), .RN(n5963), .Q(n383)
         );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n3712), .CK(CLK), .RN(n5963), .Q(n382)
         );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n3713), .CK(CLK), .RN(n5963), .Q(n381)
         );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n3714), .CK(CLK), .RN(n5963), .Q(n380)
         );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n3715), .CK(CLK), .RN(n5963), .Q(n379)
         );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n3716), .CK(CLK), .RN(n5963), .Q(n378)
         );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n3717), .CK(CLK), .RN(n5962), .Q(n377)
         );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n3718), .CK(CLK), .RN(n5962), .Q(n376)
         );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n3719), .CK(CLK), .RN(n5962), .Q(n375)
         );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n3720), .CK(CLK), .RN(n5962), .Q(n374)
         );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n3721), .CK(CLK), .RN(n5962), .Q(n373)
         );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n3722), .CK(CLK), .RN(n5962), .Q(n372)
         );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n3723), .CK(CLK), .RN(n5962), .Q(n371)
         );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n3724), .CK(CLK), .RN(n5962), .Q(n370)
         );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n3725), .CK(CLK), .RN(n5962), .Q(n369)
         );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n3726), .CK(CLK), .RN(n5962), .Q(n368)
         );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n3727), .CK(CLK), .RN(n5962), .Q(n367)
         );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n3728), .CK(CLK), .RN(n5961), .Q(n366)
         );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n3729), .CK(CLK), .RN(n5961), .Q(n365)
         );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n3730), .CK(CLK), .RN(n5961), .Q(n364)
         );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n3731), .CK(CLK), .RN(n5961), .Q(n363)
         );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n3732), .CK(CLK), .RN(n5961), .Q(n362)
         );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n3733), .CK(CLK), .RN(n5961), .Q(n361)
         );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n3734), .CK(CLK), .RN(n5961), .Q(n360)
         );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n3735), .CK(CLK), .RN(n5961), .Q(n359)
         );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n3736), .CK(CLK), .RN(n5961), .Q(n358)
         );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n3737), .CK(CLK), .RN(n5961), .Q(n357)
         );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n3738), .CK(CLK), .RN(n5961), .Q(n356)
         );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n3739), .CK(CLK), .RN(n5960), .Q(n355)
         );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n3740), .CK(CLK), .RN(n5960), .Q(n354)
         );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n3741), .CK(CLK), .RN(n5960), .Q(n353)
         );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n3742), .CK(CLK), .RN(n5960), .Q(n352)
         );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n3743), .CK(CLK), .RN(n5960), .Q(n351)
         );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n3744), .CK(CLK), .RN(n5960), .Q(n350)
         );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n3745), .CK(CLK), .RN(n5960), .Q(n349)
         );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n3746), .CK(CLK), .RN(n5960), .Q(n348)
         );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n3747), .CK(CLK), .RN(n5960), .Q(n347)
         );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n3748), .CK(CLK), .RN(n5960), .Q(n346)
         );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n3749), .CK(CLK), .RN(n5960), .Q(n345)
         );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n3750), .CK(CLK), .RN(n5959), .Q(n344)
         );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n3751), .CK(CLK), .RN(n5959), .Q(n343)
         );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n3752), .CK(CLK), .RN(n5959), .Q(n342)
         );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n3753), .CK(CLK), .RN(n5959), .Q(n341)
         );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n3754), .CK(CLK), .RN(n5959), .Q(n340)
         );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n3755), .CK(CLK), .RN(n5959), .Q(n339)
         );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n3756), .CK(CLK), .RN(n5959), .Q(n338)
         );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n3757), .CK(CLK), .RN(n5959), .Q(n337)
         );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n3758), .CK(CLK), .RN(n5959), .Q(n336)
         );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n3759), .CK(CLK), .RN(n5959), .Q(n335)
         );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n3760), .CK(CLK), .RN(n5959), .Q(n334)
         );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n3761), .CK(CLK), .RN(n5958), .Q(n333)
         );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n3762), .CK(CLK), .RN(n5958), .Q(n332)
         );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n3763), .CK(CLK), .RN(n5958), .Q(n331)
         );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n3764), .CK(CLK), .RN(n5958), .Q(n330)
         );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n3765), .CK(CLK), .RN(n5958), .Q(n329)
         );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n3766), .CK(CLK), .RN(n5958), .Q(n328)
         );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n3767), .CK(CLK), .RN(n5958), .Q(n327)
         );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n3768), .CK(CLK), .RN(n5958), .Q(n326)
         );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n3769), .CK(CLK), .RN(n5958), .Q(n325)
         );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n3770), .CK(CLK), .RN(n5958), .Q(n324)
         );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n3771), .CK(CLK), .RN(n5958), .Q(n323)
         );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n3772), .CK(CLK), .RN(n5957), .Q(n322)
         );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n3773), .CK(CLK), .RN(n5957), .Q(n321)
         );
  DFFR_X1 \OUT1_reg[31]  ( .D(n3229), .CK(CLK), .RN(n5957), .Q(OUT1[31]) );
  DFFR_X1 \OUT1_reg[30]  ( .D(n3228), .CK(CLK), .RN(n5957), .Q(OUT1[30]) );
  DFFR_X1 \OUT1_reg[29]  ( .D(n3227), .CK(CLK), .RN(n5957), .Q(OUT1[29]) );
  DFFR_X1 \OUT1_reg[28]  ( .D(n3226), .CK(CLK), .RN(n5957), .Q(OUT1[28]) );
  DFFR_X1 \OUT1_reg[27]  ( .D(n3225), .CK(CLK), .RN(n5957), .Q(OUT1[27]) );
  DFFR_X1 \OUT1_reg[26]  ( .D(n3224), .CK(CLK), .RN(n5957), .Q(OUT1[26]) );
  DFFR_X1 \OUT1_reg[25]  ( .D(n3223), .CK(CLK), .RN(n5957), .Q(OUT1[25]) );
  DFFR_X1 \OUT1_reg[24]  ( .D(n3222), .CK(CLK), .RN(n5957), .Q(OUT1[24]) );
  DFFR_X1 \OUT1_reg[23]  ( .D(n3221), .CK(CLK), .RN(n5957), .Q(OUT1[23]) );
  DFFR_X1 \OUT1_reg[22]  ( .D(n3220), .CK(CLK), .RN(n5956), .Q(OUT1[22]) );
  DFFR_X1 \OUT1_reg[21]  ( .D(n3219), .CK(CLK), .RN(n5956), .Q(OUT1[21]) );
  DFFR_X1 \OUT1_reg[20]  ( .D(n3218), .CK(CLK), .RN(n5956), .Q(OUT1[20]) );
  DFFR_X1 \OUT1_reg[19]  ( .D(n3217), .CK(CLK), .RN(n5956), .Q(OUT1[19]) );
  DFFR_X1 \OUT1_reg[18]  ( .D(n3216), .CK(CLK), .RN(n5956), .Q(OUT1[18]) );
  DFFR_X1 \OUT1_reg[17]  ( .D(n3215), .CK(CLK), .RN(n5956), .Q(OUT1[17]) );
  DFFR_X1 \OUT1_reg[16]  ( .D(n3214), .CK(CLK), .RN(n5956), .Q(OUT1[16]) );
  DFFR_X1 \OUT1_reg[15]  ( .D(n3213), .CK(CLK), .RN(n5956), .Q(OUT1[15]) );
  DFFR_X1 \OUT1_reg[14]  ( .D(n3212), .CK(CLK), .RN(n5956), .Q(OUT1[14]) );
  DFFR_X1 \OUT1_reg[13]  ( .D(n3211), .CK(CLK), .RN(n5956), .Q(OUT1[13]) );
  DFFR_X1 \OUT1_reg[12]  ( .D(n3210), .CK(CLK), .RN(n5956), .Q(OUT1[12]) );
  DFFR_X1 \OUT1_reg[11]  ( .D(n3209), .CK(CLK), .RN(n5955), .Q(OUT1[11]) );
  DFFR_X1 \OUT1_reg[10]  ( .D(n3208), .CK(CLK), .RN(n5955), .Q(OUT1[10]) );
  DFFR_X1 \OUT1_reg[9]  ( .D(n3207), .CK(CLK), .RN(n5955), .Q(OUT1[9]) );
  DFFR_X1 \OUT1_reg[8]  ( .D(n3206), .CK(CLK), .RN(n5955), .Q(OUT1[8]) );
  DFFR_X1 \OUT1_reg[7]  ( .D(n3205), .CK(CLK), .RN(n5955), .Q(OUT1[7]) );
  DFFR_X1 \OUT1_reg[6]  ( .D(n3204), .CK(CLK), .RN(n5955), .Q(OUT1[6]) );
  DFFR_X1 \OUT1_reg[5]  ( .D(n3203), .CK(CLK), .RN(n5955), .Q(OUT1[5]) );
  DFFR_X1 \OUT1_reg[4]  ( .D(n3202), .CK(CLK), .RN(n5955), .Q(OUT1[4]) );
  DFFR_X1 \OUT1_reg[3]  ( .D(n3201), .CK(CLK), .RN(n5955), .Q(OUT1[3]) );
  DFFR_X1 \OUT1_reg[2]  ( .D(n3200), .CK(CLK), .RN(n5955), .Q(OUT1[2]) );
  DFFR_X1 \OUT1_reg[1]  ( .D(n3199), .CK(CLK), .RN(n5955), .Q(OUT1[1]) );
  DFFR_X1 \OUT1_reg[0]  ( .D(n3198), .CK(CLK), .RN(n5954), .Q(OUT1[0]) );
  DFFR_X1 \OUT2_reg[31]  ( .D(n3197), .CK(CLK), .RN(n5954), .Q(OUT2[31]) );
  DFFR_X1 \OUT2_reg[30]  ( .D(n3196), .CK(CLK), .RN(n5954), .Q(OUT2[30]) );
  DFFR_X1 \OUT2_reg[29]  ( .D(n3195), .CK(CLK), .RN(n5954), .Q(OUT2[29]) );
  DFFR_X1 \OUT2_reg[28]  ( .D(n3194), .CK(CLK), .RN(n5954), .Q(OUT2[28]) );
  DFFR_X1 \OUT2_reg[27]  ( .D(n3193), .CK(CLK), .RN(n5954), .Q(OUT2[27]) );
  DFFR_X1 \OUT2_reg[26]  ( .D(n3192), .CK(CLK), .RN(n5954), .Q(OUT2[26]) );
  DFFR_X1 \OUT2_reg[25]  ( .D(n3191), .CK(CLK), .RN(n5954), .Q(OUT2[25]) );
  DFFR_X1 \OUT2_reg[24]  ( .D(n3190), .CK(CLK), .RN(n5954), .Q(OUT2[24]) );
  DFFR_X1 \OUT2_reg[23]  ( .D(n3189), .CK(CLK), .RN(n5954), .Q(OUT2[23]) );
  DFFR_X1 \OUT2_reg[22]  ( .D(n3188), .CK(CLK), .RN(n5954), .Q(OUT2[22]) );
  DFFR_X1 \OUT2_reg[21]  ( .D(n3187), .CK(CLK), .RN(n5953), .Q(OUT2[21]) );
  DFFR_X1 \OUT2_reg[20]  ( .D(n3186), .CK(CLK), .RN(n5953), .Q(OUT2[20]) );
  DFFR_X1 \OUT2_reg[19]  ( .D(n3185), .CK(CLK), .RN(n5953), .Q(OUT2[19]) );
  DFFR_X1 \OUT2_reg[18]  ( .D(n3184), .CK(CLK), .RN(n5953), .Q(OUT2[18]) );
  DFFR_X1 \OUT2_reg[17]  ( .D(n3183), .CK(CLK), .RN(n5953), .Q(OUT2[17]) );
  DFFR_X1 \OUT2_reg[16]  ( .D(n3182), .CK(CLK), .RN(n5953), .Q(OUT2[16]) );
  DFFR_X1 \OUT2_reg[15]  ( .D(n3181), .CK(CLK), .RN(n5953), .Q(OUT2[15]) );
  DFFR_X1 \OUT2_reg[14]  ( .D(n3180), .CK(CLK), .RN(n5953), .Q(OUT2[14]) );
  DFFR_X1 \OUT2_reg[13]  ( .D(n3179), .CK(CLK), .RN(n5953), .Q(OUT2[13]) );
  DFFR_X1 \OUT2_reg[12]  ( .D(n3178), .CK(CLK), .RN(n5953), .Q(OUT2[12]) );
  DFFR_X1 \OUT2_reg[11]  ( .D(n3177), .CK(CLK), .RN(n5953), .Q(OUT2[11]) );
  DFFR_X1 \OUT2_reg[10]  ( .D(n3176), .CK(CLK), .RN(n5952), .Q(OUT2[10]) );
  DFFR_X1 \OUT2_reg[9]  ( .D(n3175), .CK(CLK), .RN(n5952), .Q(OUT2[9]) );
  DFFR_X1 \OUT2_reg[8]  ( .D(n3174), .CK(CLK), .RN(n5952), .Q(OUT2[8]) );
  DFFR_X1 \OUT2_reg[7]  ( .D(n3173), .CK(CLK), .RN(n5952), .Q(OUT2[7]) );
  DFFR_X1 \OUT2_reg[6]  ( .D(n3172), .CK(CLK), .RN(n5952), .Q(OUT2[6]) );
  DFFR_X1 \OUT2_reg[5]  ( .D(n3171), .CK(CLK), .RN(n5952), .Q(OUT2[5]) );
  DFFR_X1 \OUT2_reg[4]  ( .D(n3170), .CK(CLK), .RN(n5952), .Q(OUT2[4]) );
  DFFR_X1 \OUT2_reg[3]  ( .D(n3169), .CK(CLK), .RN(n5952), .Q(OUT2[3]) );
  DFFR_X1 \OUT2_reg[2]  ( .D(n3168), .CK(CLK), .RN(n5952), .Q(OUT2[2]) );
  DFFR_X1 \OUT2_reg[1]  ( .D(n3167), .CK(CLK), .RN(n5952), .Q(OUT2[1]) );
  DFFR_X1 \OUT2_reg[0]  ( .D(n3166), .CK(CLK), .RN(n5952), .Q(OUT2[0]) );
  NOR2_X1 U4 ( .A1(n6621), .A2(n6622), .ZN(n5332) );
  OR3_X1 U5 ( .A1(n5293), .A2(n5290), .A3(n5292), .ZN(n6621) );
  OR3_X1 U7 ( .A1(n5289), .A2(n6620), .A3(n5288), .ZN(n6622) );
  NOR2_X1 U8 ( .A1(n6623), .A2(n6624), .ZN(n4430) );
  OR3_X1 U9 ( .A1(n4391), .A2(n4388), .A3(n4390), .ZN(n6623) );
  OR3_X1 U10 ( .A1(n4387), .A2(n6620), .A3(n4386), .ZN(n6624) );
  AND2_X1 U11 ( .A1(n2307), .A2(ADD_WR[1]), .ZN(n1658) );
  AND2_X1 U12 ( .A1(n2341), .A2(ADD_WR[1]), .ZN(n1624) );
  AND2_X1 U13 ( .A1(n5353), .A2(ADD_WR[1]), .ZN(n1590) );
  AND2_X1 U14 ( .A1(n2419), .A2(ADD_WR[1]), .ZN(n1555) );
  NAND4_X1 U15 ( .A1(n5300), .A2(n5301), .A3(n5302), .A4(n5303), .ZN(n5276) );
  NAND4_X1 U16 ( .A1(n5258), .A2(n5259), .A3(n5260), .A4(n5261), .ZN(n5250) );
  NAND4_X1 U17 ( .A1(n5232), .A2(n5233), .A3(n5234), .A4(n5235), .ZN(n5224) );
  NAND4_X1 U19 ( .A1(n5206), .A2(n5207), .A3(n5208), .A4(n5209), .ZN(n5198) );
  NAND4_X1 U21 ( .A1(n5180), .A2(n5181), .A3(n5182), .A4(n5183), .ZN(n5172) );
  NAND4_X1 U22 ( .A1(n5154), .A2(n5155), .A3(n5156), .A4(n5157), .ZN(n5146) );
  NAND4_X1 U23 ( .A1(n5128), .A2(n5129), .A3(n5130), .A4(n5131), .ZN(n5120) );
  NAND4_X1 U24 ( .A1(n5102), .A2(n5103), .A3(n5104), .A4(n5105), .ZN(n5094) );
  NAND4_X1 U25 ( .A1(n5076), .A2(n5077), .A3(n5078), .A4(n5079), .ZN(n5068) );
  NAND4_X1 U26 ( .A1(n5050), .A2(n5051), .A3(n5052), .A4(n5053), .ZN(n5042) );
  NAND4_X1 U27 ( .A1(n5024), .A2(n5025), .A3(n5026), .A4(n5027), .ZN(n5016) );
  NAND4_X1 U29 ( .A1(n4998), .A2(n4999), .A3(n5000), .A4(n5001), .ZN(n4990) );
  NAND4_X1 U30 ( .A1(n4972), .A2(n4973), .A3(n4974), .A4(n4975), .ZN(n4964) );
  NAND4_X1 U31 ( .A1(n4946), .A2(n4947), .A3(n4948), .A4(n4949), .ZN(n4938) );
  NAND4_X1 U32 ( .A1(n4920), .A2(n4921), .A3(n4922), .A4(n4923), .ZN(n4912) );
  NAND4_X1 U33 ( .A1(n4894), .A2(n4895), .A3(n4896), .A4(n4897), .ZN(n4886) );
  NAND4_X1 U34 ( .A1(n4868), .A2(n4869), .A3(n4870), .A4(n4871), .ZN(n4860) );
  NAND4_X1 U35 ( .A1(n4842), .A2(n4843), .A3(n4844), .A4(n4845), .ZN(n4834) );
  NAND4_X1 U36 ( .A1(n4816), .A2(n4817), .A3(n4818), .A4(n4819), .ZN(n4808) );
  NAND4_X1 U37 ( .A1(n4790), .A2(n4791), .A3(n4792), .A4(n4793), .ZN(n4782) );
  NAND4_X1 U38 ( .A1(n4764), .A2(n4765), .A3(n4766), .A4(n4767), .ZN(n4756) );
  NAND4_X1 U39 ( .A1(n4738), .A2(n4739), .A3(n4740), .A4(n4741), .ZN(n4730) );
  NAND4_X1 U40 ( .A1(n4712), .A2(n4713), .A3(n4714), .A4(n4715), .ZN(n4704) );
  NAND4_X1 U41 ( .A1(n4686), .A2(n4687), .A3(n4688), .A4(n4689), .ZN(n4678) );
  NAND4_X1 U42 ( .A1(n4660), .A2(n4661), .A3(n4662), .A4(n4663), .ZN(n4652) );
  NAND4_X1 U43 ( .A1(n4634), .A2(n4635), .A3(n4636), .A4(n4637), .ZN(n4626) );
  NAND4_X1 U45 ( .A1(n4608), .A2(n4609), .A3(n4610), .A4(n4611), .ZN(n4600) );
  NAND4_X1 U47 ( .A1(n4582), .A2(n4583), .A3(n4584), .A4(n4585), .ZN(n4574) );
  NAND4_X1 U48 ( .A1(n4556), .A2(n4557), .A3(n4558), .A4(n4559), .ZN(n4548) );
  NAND4_X1 U49 ( .A1(n4530), .A2(n4531), .A3(n4532), .A4(n4533), .ZN(n4522) );
  NAND4_X1 U51 ( .A1(n4504), .A2(n4505), .A3(n4506), .A4(n4507), .ZN(n4496) );
  NAND4_X1 U52 ( .A1(n4455), .A2(n4456), .A3(n4457), .A4(n4458), .ZN(n4438) );
  NAND4_X1 U55 ( .A1(n4398), .A2(n4399), .A3(n4400), .A4(n4401), .ZN(n4374) );
  NAND4_X1 U56 ( .A1(n4356), .A2(n4357), .A3(n4358), .A4(n4359), .ZN(n4348) );
  NAND4_X1 U57 ( .A1(n4330), .A2(n4331), .A3(n4332), .A4(n4333), .ZN(n4322) );
  NAND4_X1 U61 ( .A1(n4304), .A2(n4305), .A3(n4306), .A4(n4307), .ZN(n4296) );
  NAND4_X1 U62 ( .A1(n4278), .A2(n4279), .A3(n4280), .A4(n4281), .ZN(n4270) );
  NAND4_X1 U63 ( .A1(n4252), .A2(n4253), .A3(n4254), .A4(n4255), .ZN(n4244) );
  NAND4_X1 U64 ( .A1(n4226), .A2(n4227), .A3(n4228), .A4(n4229), .ZN(n4218) );
  NAND4_X1 U65 ( .A1(n4200), .A2(n4201), .A3(n4202), .A4(n4203), .ZN(n4192) );
  NAND4_X1 U66 ( .A1(n3982), .A2(n3983), .A3(n3984), .A4(n3985), .ZN(n3974) );
  NAND4_X1 U69 ( .A1(n3956), .A2(n3957), .A3(n3958), .A4(n3959), .ZN(n3948) );
  NAND4_X1 U71 ( .A1(n3930), .A2(n3931), .A3(n3932), .A4(n3933), .ZN(n3922) );
  NAND4_X1 U72 ( .A1(n3040), .A2(n3041), .A3(n3042), .A4(n3043), .ZN(n3032) );
  NAND4_X1 U73 ( .A1(n3014), .A2(n3015), .A3(n3016), .A4(n3017), .ZN(n3006) );
  NAND4_X1 U74 ( .A1(n2988), .A2(n2989), .A3(n2990), .A4(n2991), .ZN(n2980) );
  NAND4_X1 U75 ( .A1(n2962), .A2(n2963), .A3(n2964), .A4(n2965), .ZN(n2954) );
  NAND4_X1 U77 ( .A1(n2936), .A2(n2937), .A3(n2938), .A4(n2939), .ZN(n2928) );
  NAND4_X1 U78 ( .A1(n2910), .A2(n2911), .A3(n2912), .A4(n2913), .ZN(n2902) );
  NAND4_X1 U79 ( .A1(n2884), .A2(n2885), .A3(n2886), .A4(n2887), .ZN(n2876) );
  NAND4_X1 U80 ( .A1(n2858), .A2(n2859), .A3(n2860), .A4(n2861), .ZN(n2850) );
  NAND4_X1 U82 ( .A1(n2832), .A2(n2833), .A3(n2834), .A4(n2835), .ZN(n2800) );
  NAND4_X1 U83 ( .A1(n2782), .A2(n2783), .A3(n2784), .A4(n2785), .ZN(n2774) );
  NAND4_X1 U84 ( .A1(n2756), .A2(n2757), .A3(n2758), .A4(n2759), .ZN(n2748) );
  NAND4_X1 U85 ( .A1(n2730), .A2(n2731), .A3(n2732), .A4(n2733), .ZN(n2722) );
  NAND4_X1 U86 ( .A1(n2704), .A2(n2705), .A3(n2706), .A4(n2707), .ZN(n2696) );
  NAND4_X1 U87 ( .A1(n2678), .A2(n2679), .A3(n2680), .A4(n2681), .ZN(n2670) );
  NAND4_X1 U89 ( .A1(n2652), .A2(n2653), .A3(n2654), .A4(n2655), .ZN(n2644) );
  NAND4_X1 U90 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(n2618) );
  NAND4_X1 U91 ( .A1(n2600), .A2(n2601), .A3(n2602), .A4(n2603), .ZN(n2592) );
  NAND4_X1 U92 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2577), .ZN(n2566) );
  NAND4_X1 U93 ( .A1(n2548), .A2(n2549), .A3(n2550), .A4(n2551), .ZN(n2540) );
  NAND4_X1 U94 ( .A1(n2522), .A2(n2523), .A3(n2524), .A4(n2525), .ZN(n2514) );
  NAND4_X1 U95 ( .A1(n2473), .A2(n2474), .A3(n2475), .A4(n2476), .ZN(n2456) );
endmodule


module sign_ext_N_IN026_N_IN116_N_OUT32 ( ctrl_in, zero_padding, data_in, 
        data_ext );
  input [25:0] data_in;
  output [31:0] data_ext;
  input ctrl_in, zero_padding;
  wire   \data_ext[31] , \data_in[15] , \data_in[14] , \data_in[13] ,
         \data_in[12] , \data_in[11] , \data_in[10] , \data_in[9] ,
         \data_in[8] , \data_in[7] , \data_in[6] , \data_in[5] , \data_in[4] ,
         \data_in[3] , \data_in[2] , \data_in[1] , \data_in[0] , n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  assign data_ext[25] = \data_ext[31] ;
  assign data_ext[26] = \data_ext[31] ;
  assign data_ext[27] = \data_ext[31] ;
  assign data_ext[28] = \data_ext[31] ;
  assign data_ext[29] = \data_ext[31] ;
  assign data_ext[30] = \data_ext[31] ;
  assign data_ext[31] = \data_ext[31] ;
  assign data_ext[15] = \data_in[15] ;
  assign \data_in[15]  = data_in[15];
  assign data_ext[14] = \data_in[14] ;
  assign \data_in[14]  = data_in[14];
  assign data_ext[13] = \data_in[13] ;
  assign \data_in[13]  = data_in[13];
  assign data_ext[12] = \data_in[12] ;
  assign \data_in[12]  = data_in[12];
  assign data_ext[11] = \data_in[11] ;
  assign \data_in[11]  = data_in[11];
  assign data_ext[10] = \data_in[10] ;
  assign \data_in[10]  = data_in[10];
  assign data_ext[9] = \data_in[9] ;
  assign \data_in[9]  = data_in[9];
  assign data_ext[8] = \data_in[8] ;
  assign \data_in[8]  = data_in[8];
  assign data_ext[7] = \data_in[7] ;
  assign \data_in[7]  = data_in[7];
  assign data_ext[6] = \data_in[6] ;
  assign \data_in[6]  = data_in[6];
  assign data_ext[5] = \data_in[5] ;
  assign \data_in[5]  = data_in[5];
  assign data_ext[4] = \data_in[4] ;
  assign \data_in[4]  = data_in[4];
  assign data_ext[3] = \data_in[3] ;
  assign \data_in[3]  = data_in[3];
  assign data_ext[2] = \data_in[2] ;
  assign \data_in[2]  = data_in[2];
  assign data_ext[1] = \data_in[1] ;
  assign \data_in[1]  = data_in[1];
  assign data_ext[0] = \data_in[0] ;
  assign \data_in[0]  = data_in[0];

  NAND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(\data_ext[31] ) );
  NAND2_X1 U4 ( .A1(data_in[25]), .A2(n14), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n2), .A2(n4), .ZN(data_ext[24]) );
  NAND2_X1 U6 ( .A1(data_in[24]), .A2(n14), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n2), .A2(n5), .ZN(data_ext[23]) );
  NAND2_X1 U8 ( .A1(data_in[23]), .A2(n14), .ZN(n5) );
  NAND2_X1 U9 ( .A1(n2), .A2(n6), .ZN(data_ext[22]) );
  NAND2_X1 U10 ( .A1(data_in[22]), .A2(n14), .ZN(n6) );
  NAND2_X1 U11 ( .A1(n2), .A2(n7), .ZN(data_ext[21]) );
  NAND2_X1 U12 ( .A1(data_in[21]), .A2(n14), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n2), .A2(n8), .ZN(data_ext[20]) );
  NAND2_X1 U14 ( .A1(data_in[20]), .A2(n14), .ZN(n8) );
  NAND2_X1 U15 ( .A1(n2), .A2(n9), .ZN(data_ext[19]) );
  NAND2_X1 U16 ( .A1(data_in[19]), .A2(n14), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n2), .A2(n10), .ZN(data_ext[18]) );
  NAND2_X1 U18 ( .A1(data_in[18]), .A2(n14), .ZN(n10) );
  NAND2_X1 U19 ( .A1(n2), .A2(n11), .ZN(data_ext[17]) );
  NAND2_X1 U20 ( .A1(data_in[17]), .A2(n14), .ZN(n11) );
  NAND2_X1 U21 ( .A1(n2), .A2(n12), .ZN(data_ext[16]) );
  NAND2_X1 U22 ( .A1(data_in[16]), .A2(n14), .ZN(n12) );
  NAND2_X1 U23 ( .A1(n13), .A2(\data_in[15] ), .ZN(n2) );
  NOR2_X1 U24 ( .A1(zero_padding), .A2(n14), .ZN(n13) );
  INV_X1 U2 ( .A(ctrl_in), .ZN(n14) );
endmodule


module gen_mux21_N5 ( sel, x, y, m );
  input [4:0] x;
  input [4:0] y;
  output [4:0] m;
  input sel;
  wire   n7, n8, n9, n10, n11, n16;

  AOI22_X1 U7 ( .A1(x[4]), .A2(n16), .B1(y[4]), .B2(sel), .ZN(n7) );
  AOI22_X1 U8 ( .A1(x[3]), .A2(n16), .B1(y[3]), .B2(sel), .ZN(n8) );
  AOI22_X1 U9 ( .A1(x[2]), .A2(n16), .B1(y[2]), .B2(sel), .ZN(n9) );
  AOI22_X1 U10 ( .A1(x[1]), .A2(n16), .B1(y[1]), .B2(sel), .ZN(n10) );
  AOI22_X1 U11 ( .A1(x[0]), .A2(n16), .B1(y[0]), .B2(sel), .ZN(n11) );
  INV_X1 U1 ( .A(n11), .ZN(m[0]) );
  INV_X1 U2 ( .A(n10), .ZN(m[1]) );
  INV_X1 U3 ( .A(n9), .ZN(m[2]) );
  INV_X1 U4 ( .A(n8), .ZN(m[3]) );
  INV_X1 U5 ( .A(n7), .ZN(m[4]) );
  INV_X1 U6 ( .A(sel), .ZN(n16) );
endmodule



    module ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 ( 
        CLK, RST, JAL_REG31, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, WR_EN, 
        ZERO_PADDING2, I_CODE, NPC1_IN, DATA_IN, WR_ADDR_IN, REGA_OUT, 
        REGB_OUT, REGIMM_OUT, WR_ADDR_OUT, NPC1_OUT );
  input [31:0] I_CODE;
  input [31:0] NPC1_IN;
  input [31:0] DATA_IN;
  input [4:0] WR_ADDR_IN;
  output [31:0] REGA_OUT;
  output [31:0] REGB_OUT;
  output [31:0] REGIMM_OUT;
  output [4:0] WR_ADDR_OUT;
  output [31:0] NPC1_OUT;
  input CLK, RST, JAL_REG31, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, WR_EN,
         ZERO_PADDING2;

  wire   [31:0] SIGN_EXT_OUT;
  wire   [4:0] MUX_OUT;
  wire   [4:0] ADD_WR;

  OR2_X1 U1 ( .A1(JAL_REG31), .A2(WR_ADDR_IN[4]), .ZN(ADD_WR[4]) );
  OR2_X1 U2 ( .A1(JAL_REG31), .A2(WR_ADDR_IN[3]), .ZN(ADD_WR[3]) );
  OR2_X1 U3 ( .A1(JAL_REG31), .A2(WR_ADDR_IN[2]), .ZN(ADD_WR[2]) );
  OR2_X1 U4 ( .A1(JAL_REG31), .A2(WR_ADDR_IN[1]), .ZN(ADD_WR[1]) );
  OR2_X1 U5 ( .A1(JAL_REG31), .A2(WR_ADDR_IN[0]), .ZN(ADD_WR[0]) );
  gen_reg_N32_7 NPC1 ( .clk(CLK), .rst(RST), .ld(DEC_OUTREG_EN), .data_in(
        NPC1_IN), .data_out(NPC1_OUT) );
  gen_reg_N32_6 IMM ( .clk(CLK), .rst(RST), .ld(DEC_OUTREG_EN), .data_in(
        SIGN_EXT_OUT), .data_out(REGIMM_OUT) );
  gen_reg_N5_0 WR_ADDR ( .clk(CLK), .rst(RST), .ld(DEC_OUTREG_EN), .data_in(
        MUX_OUT), .data_out(WR_ADDR_OUT) );
  reg_file_Dbits32_Abits5 RF ( .CLK(CLK), .RESET(RST), .ENABLE(DEC_OUTREG_EN), 
        .RD1(RD1_EN), .RD2(RD2_EN), .WR(WR_EN), .ADD_WR(ADD_WR), .ADD_RD1(
        I_CODE[25:21]), .ADD_RD2(I_CODE[20:16]), .DATAIN(DATA_IN), .OUT1(
        REGA_OUT), .OUT2(REGB_OUT) );
  sign_ext_N_IN026_N_IN116_N_OUT32 SIGN_EXTEND ( .ctrl_in(IS_I_TYPE), 
        .zero_padding(ZERO_PADDING2), .data_in(I_CODE[25:0]), .data_ext(
        SIGN_EXT_OUT) );
  gen_mux21_N5 MUX_WR_ADDR ( .sel(IS_I_TYPE), .x(I_CODE[15:11]), .y(
        I_CODE[20:16]), .m(MUX_OUT) );
endmodule


module gen_reg_N32_5 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n99, n100, n110, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181;

  OAI21_X1 U2 ( .B1(n173), .B2(n110), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n110), .A2(data_in[23]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n174), .B2(n99), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[24]), .A2(ld), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n175), .B2(n100), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[25]), .A2(ld), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n176), .B2(n100), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[26]), .A2(n100), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n177), .B2(n110), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[27]), .A2(n100), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n178), .B2(n100), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[28]), .A2(n110), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n110), .A(n143), .ZN(n32) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n110), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n110), .A(n142), .ZN(n31) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n99), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n110), .A(n141), .ZN(n30) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n100), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n179), .B2(n110), .A(n140), .ZN(n3) );
  NAND2_X1 U21 ( .A1(data_in[29]), .A2(n110), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n153), .B2(n99), .A(n139), .ZN(n29) );
  NAND2_X1 U23 ( .A1(data_in[3]), .A2(n100), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n154), .B2(n110), .A(n138), .ZN(n28) );
  NAND2_X1 U25 ( .A1(data_in[4]), .A2(n99), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n155), .B2(n100), .A(n137), .ZN(n27) );
  NAND2_X1 U27 ( .A1(data_in[5]), .A2(n100), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n156), .B2(n99), .A(n136), .ZN(n26) );
  NAND2_X1 U29 ( .A1(data_in[6]), .A2(n99), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n157), .B2(n110), .A(n135), .ZN(n25) );
  NAND2_X1 U31 ( .A1(data_in[7]), .A2(n100), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n158), .B2(n110), .A(n134), .ZN(n24) );
  NAND2_X1 U33 ( .A1(data_in[8]), .A2(n99), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n159), .B2(n99), .A(n133), .ZN(n23) );
  NAND2_X1 U35 ( .A1(data_in[9]), .A2(n100), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n160), .B2(n110), .A(n132), .ZN(n22) );
  NAND2_X1 U37 ( .A1(data_in[10]), .A2(n99), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n161), .B2(n110), .A(n131), .ZN(n21) );
  NAND2_X1 U39 ( .A1(data_in[11]), .A2(n100), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n162), .B2(n110), .A(n130), .ZN(n20) );
  NAND2_X1 U41 ( .A1(data_in[12]), .A2(n99), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n180), .B2(n99), .A(n129), .ZN(n2) );
  NAND2_X1 U43 ( .A1(data_in[30]), .A2(n110), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n163), .B2(n100), .A(n128), .ZN(n19) );
  NAND2_X1 U45 ( .A1(data_in[13]), .A2(n100), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n164), .B2(n100), .A(n127), .ZN(n18) );
  NAND2_X1 U47 ( .A1(data_in[14]), .A2(n110), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n165), .B2(n99), .A(n126), .ZN(n17) );
  NAND2_X1 U49 ( .A1(data_in[15]), .A2(n100), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n166), .B2(n99), .A(n125), .ZN(n16) );
  NAND2_X1 U51 ( .A1(data_in[16]), .A2(n99), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n167), .B2(n100), .A(n124), .ZN(n15) );
  NAND2_X1 U53 ( .A1(data_in[17]), .A2(ld), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n168), .B2(n110), .A(n123), .ZN(n14) );
  NAND2_X1 U55 ( .A1(data_in[18]), .A2(n99), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n169), .B2(n100), .A(n122), .ZN(n13) );
  NAND2_X1 U57 ( .A1(data_in[19]), .A2(n110), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n170), .B2(n110), .A(n121), .ZN(n12) );
  NAND2_X1 U59 ( .A1(data_in[20]), .A2(n110), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n171), .B2(n99), .A(n120), .ZN(n11) );
  NAND2_X1 U61 ( .A1(data_in[21]), .A2(n99), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n172), .B2(n110), .A(n119), .ZN(n10) );
  NAND2_X1 U63 ( .A1(data_in[22]), .A2(n100), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n181), .B2(n99), .A(n118), .ZN(n1) );
  NAND2_X1 U65 ( .A1(data_in[31]), .A2(n99), .ZN(n118) );
  CLKBUF_X1 U67 ( .A(n110), .Z(n99) );
  CLKBUF_X1 U71 ( .A(n110), .Z(n100) );
  CLKBUF_X1 U82 ( .A(ld), .Z(n110) );
  DFFR_X1 \data_out_reg[31]  ( .D(n1), .CK(clk), .RN(rst), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n2), .CK(clk), .RN(rst), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n3), .CK(clk), .RN(rst), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n6), .CK(clk), .RN(rst), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n7), .CK(clk), .RN(rst), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n8), .CK(clk), .RN(rst), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n9), .CK(clk), .RN(rst), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n10), .CK(clk), .RN(rst), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n11), .CK(clk), .RN(rst), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n12), .CK(clk), .RN(rst), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n13), .CK(clk), .RN(rst), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n14), .CK(clk), .RN(rst), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n15), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n16), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n17), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n23), .CK(clk), .RN(rst), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n24), .CK(clk), .RN(rst), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n25), .CK(clk), .RN(rst), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n26), .CK(clk), .RN(rst), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n27), .CK(clk), .RN(rst), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n28), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n29), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n30), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n31), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module zero_check_N32 ( data_in, ctrl_out );
  input [31:0] data_in;
  output ctrl_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  NOR4_X1 U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(ctrl_out) );
  NAND2_X1 U2 ( .A1(n5), .A2(n6), .ZN(n4) );
  NOR4_X1 U3 ( .A1(data_in[16]), .A2(data_in[15]), .A3(data_in[14]), .A4(
        data_in[13]), .ZN(n6) );
  NOR4_X1 U4 ( .A1(data_in[12]), .A2(data_in[11]), .A3(data_in[10]), .A4(
        data_in[0]), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(n3) );
  NOR4_X1 U6 ( .A1(data_in[23]), .A2(data_in[22]), .A3(data_in[21]), .A4(
        data_in[20]), .ZN(n8) );
  NOR4_X1 U7 ( .A1(data_in[1]), .A2(data_in[19]), .A3(data_in[18]), .A4(
        data_in[17]), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n9), .A2(n10), .ZN(n2) );
  NOR4_X1 U9 ( .A1(data_in[30]), .A2(data_in[2]), .A3(data_in[29]), .A4(
        data_in[28]), .ZN(n10) );
  NOR4_X1 U10 ( .A1(data_in[27]), .A2(data_in[26]), .A3(data_in[25]), .A4(
        data_in[24]), .ZN(n9) );
  NAND2_X1 U11 ( .A1(n11), .A2(n12), .ZN(n1) );
  NOR4_X1 U12 ( .A1(data_in[9]), .A2(data_in[8]), .A3(data_in[7]), .A4(
        data_in[6]), .ZN(n12) );
  NOR4_X1 U13 ( .A1(data_in[5]), .A2(data_in[4]), .A3(data_in[3]), .A4(
        data_in[31]), .ZN(n11) );
endmodule


module cond_branch ( cond_in, jump_in, ctrl_in, ctrl_out );
  input cond_in, jump_in, ctrl_in;
  output ctrl_out;
  wire   n1;

  XNOR2_X1 U2 ( .A(ctrl_in), .B(cond_in), .ZN(n1) );
  AND2_X1 U1 ( .A1(n1), .A2(jump_in), .ZN(ctrl_out) );
endmodule


module gen_mux21_N32_0 ( sel, x, y, m );
  input [31:0] x;
  input [31:0] y;
  output [31:0] m;
  input sel;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, net74010, net74997, net74991, net76453, net83431,
         net83447, net83646, net88215, n54;
  assign m[1] = net74010;

  AOI22_X1 U34 ( .A1(x[9]), .A2(net76453), .B1(y[9]), .B2(net83646), .ZN(n34)
         );
  AOI22_X1 U35 ( .A1(x[8]), .A2(net76453), .B1(y[8]), .B2(net74997), .ZN(n35)
         );
  AOI22_X1 U36 ( .A1(x[7]), .A2(net76453), .B1(y[7]), .B2(net74997), .ZN(n36)
         );
  AOI22_X1 U37 ( .A1(x[6]), .A2(net76453), .B1(y[6]), .B2(net74997), .ZN(n37)
         );
  AOI22_X1 U38 ( .A1(x[5]), .A2(net76453), .B1(y[5]), .B2(net83646), .ZN(n38)
         );
  AOI22_X1 U39 ( .A1(x[4]), .A2(net76453), .B1(y[4]), .B2(net83646), .ZN(n39)
         );
  AOI22_X1 U40 ( .A1(x[3]), .A2(net74991), .B1(y[3]), .B2(net74997), .ZN(n40)
         );
  AOI22_X1 U41 ( .A1(x[31]), .A2(net76453), .B1(y[31]), .B2(net88215), .ZN(n41) );
  AOI22_X1 U42 ( .A1(x[30]), .A2(net76453), .B1(y[30]), .B2(net88215), .ZN(n42) );
  AOI22_X1 U43 ( .A1(x[2]), .A2(net74991), .B1(net83447), .B2(y[2]), .ZN(n43)
         );
  AOI22_X1 U44 ( .A1(x[29]), .A2(net76453), .B1(y[29]), .B2(net88215), .ZN(n44) );
  AOI22_X1 U45 ( .A1(x[28]), .A2(net76453), .B1(y[28]), .B2(net83646), .ZN(n45) );
  AOI22_X1 U46 ( .A1(x[27]), .A2(net76453), .B1(y[27]), .B2(net83646), .ZN(n46) );
  AOI22_X1 U47 ( .A1(x[26]), .A2(net76453), .B1(y[26]), .B2(net83646), .ZN(n47) );
  AOI22_X1 U48 ( .A1(x[25]), .A2(net76453), .B1(y[25]), .B2(net83646), .ZN(n48) );
  AOI22_X1 U49 ( .A1(x[24]), .A2(net76453), .B1(y[24]), .B2(net83646), .ZN(n49) );
  AOI22_X1 U50 ( .A1(x[23]), .A2(net76453), .B1(y[23]), .B2(net83646), .ZN(n50) );
  AOI22_X1 U51 ( .A1(x[22]), .A2(net76453), .B1(y[22]), .B2(net83646), .ZN(n51) );
  AOI22_X1 U52 ( .A1(x[21]), .A2(net76453), .B1(y[21]), .B2(net88215), .ZN(n52) );
  AOI22_X1 U53 ( .A1(x[20]), .A2(net76453), .B1(y[20]), .B2(net88215), .ZN(n53) );
  AOI22_X1 U55 ( .A1(x[19]), .A2(net76453), .B1(y[19]), .B2(net88215), .ZN(n55) );
  AOI22_X1 U56 ( .A1(x[18]), .A2(net76453), .B1(y[18]), .B2(net88215), .ZN(n56) );
  AOI22_X1 U57 ( .A1(x[17]), .A2(net76453), .B1(y[17]), .B2(net88215), .ZN(n57) );
  AOI22_X1 U58 ( .A1(x[16]), .A2(net76453), .B1(y[16]), .B2(net88215), .ZN(n58) );
  AOI22_X1 U59 ( .A1(x[15]), .A2(net76453), .B1(y[15]), .B2(net88215), .ZN(n59) );
  AOI22_X1 U60 ( .A1(x[14]), .A2(net76453), .B1(y[14]), .B2(net88215), .ZN(n60) );
  AOI22_X1 U61 ( .A1(x[13]), .A2(net76453), .B1(y[13]), .B2(net88215), .ZN(n61) );
  AOI22_X1 U62 ( .A1(x[12]), .A2(net76453), .B1(y[12]), .B2(net88215), .ZN(n62) );
  AOI22_X1 U63 ( .A1(x[11]), .A2(net76453), .B1(y[11]), .B2(net88215), .ZN(n63) );
  AOI22_X1 U64 ( .A1(x[10]), .A2(net76453), .B1(y[10]), .B2(net88215), .ZN(n64) );
  AOI22_X1 U65 ( .A1(net74991), .A2(x[0]), .B1(net83431), .B2(y[0]), .ZN(n65)
         );
  AOI22_X1 U54 ( .A1(net74991), .A2(x[1]), .B1(net83431), .B2(y[1]), .ZN(n54)
         );
  INV_X1 U2 ( .A(n54), .ZN(net74010) );
  CLKBUF_X1 U4 ( .A(net83447), .Z(net74997) );
  INV_X1 U5 ( .A(sel), .ZN(net74991) );
  CLKBUF_X1 U6 ( .A(sel), .Z(net83431) );
  CLKBUF_X1 U7 ( .A(net83447), .Z(net88215) );
  INV_X1 U15 ( .A(n40), .ZN(m[3]) );
  INV_X1 U16 ( .A(n43), .ZN(m[2]) );
  INV_X1 U19 ( .A(n35), .ZN(m[8]) );
  INV_X1 U20 ( .A(n64), .ZN(m[10]) );
  INV_X1 U21 ( .A(n63), .ZN(m[11]) );
  INV_X1 U22 ( .A(n57), .ZN(m[17]) );
  INV_X1 U23 ( .A(n59), .ZN(m[15]) );
  INV_X1 U24 ( .A(n58), .ZN(m[16]) );
  INV_X1 U25 ( .A(n61), .ZN(m[13]) );
  INV_X1 U26 ( .A(n60), .ZN(m[14]) );
  INV_X1 U27 ( .A(n37), .ZN(m[6]) );
  INV_X1 U28 ( .A(n62), .ZN(m[12]) );
  INV_X1 U29 ( .A(n39), .ZN(m[4]) );
  INV_X1 U30 ( .A(n38), .ZN(m[5]) );
  INV_X1 U31 ( .A(n55), .ZN(m[19]) );
  INV_X1 U32 ( .A(n56), .ZN(m[18]) );
  INV_X1 U33 ( .A(n53), .ZN(m[20]) );
  INV_X1 U66 ( .A(n49), .ZN(m[24]) );
  INV_X1 U67 ( .A(n50), .ZN(m[23]) );
  INV_X1 U68 ( .A(n42), .ZN(m[30]) );
  INV_X1 U69 ( .A(n44), .ZN(m[29]) );
  INV_X1 U70 ( .A(n51), .ZN(m[22]) );
  INV_X1 U71 ( .A(n47), .ZN(m[26]) );
  INV_X1 U72 ( .A(n45), .ZN(m[28]) );
  INV_X1 U73 ( .A(n46), .ZN(m[27]) );
  INV_X1 U74 ( .A(n48), .ZN(m[25]) );
  INV_X1 U75 ( .A(n41), .ZN(m[31]) );
  INV_X1 U76 ( .A(n52), .ZN(m[21]) );
  INV_X1 U77 ( .A(n65), .ZN(m[0]) );
  BUF_X1 U1 ( .A(net74997), .Z(net83646) );
  INV_X1 U3 ( .A(n34), .ZN(m[9]) );
  INV_X1 U8 ( .A(n36), .ZN(m[7]) );
  CLKBUF_X1 U9 ( .A(net83431), .Z(net83447) );
  CLKBUF_X3 U10 ( .A(net74991), .Z(net76453) );
endmodule


module gen_mux21_N32_2 ( sel, x, y, m );
  input [31:0] x;
  input [31:0] y;
  output [31:0] m;
  input sel;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n64,
         net74042, net74045, net74046, net74049, net74051, net74052, net74053,
         net74054, net74056, net75023, net82700, net82897, net83357, net83766,
         n65, net88219, net94624, net75011, net107657, n62, net112175, n63,
         net76465, net75025, net75015, n34;
  assign m[0] = net74042;
  assign m[3] = net74045;
  assign m[4] = net74046;
  assign m[7] = net74049;
  assign m[9] = net74051;
  assign m[10] = net74052;
  assign m[11] = net74053;
  assign m[12] = net74054;
  assign m[14] = net74056;

  AOI22_X1 U35 ( .A1(x[8]), .A2(net88219), .B1(y[8]), .B2(net94624), .ZN(n35)
         );
  AOI22_X1 U37 ( .A1(x[6]), .A2(net88219), .B1(y[6]), .B2(net94624), .ZN(n37)
         );
  AOI22_X1 U38 ( .A1(x[5]), .A2(net88219), .B1(net94624), .B2(y[5]), .ZN(n38)
         );
  AOI22_X1 U41 ( .A1(x[31]), .A2(net82897), .B1(y[31]), .B2(net83766), .ZN(n41) );
  AOI22_X1 U42 ( .A1(x[30]), .A2(net82897), .B1(y[30]), .B2(net83766), .ZN(n42) );
  AOI22_X1 U43 ( .A1(x[2]), .A2(net112175), .B1(y[2]), .B2(net83357), .ZN(n43)
         );
  AOI22_X1 U44 ( .A1(x[29]), .A2(net82897), .B1(y[29]), .B2(net83766), .ZN(n44) );
  AOI22_X1 U45 ( .A1(x[28]), .A2(net82897), .B1(y[28]), .B2(net83766), .ZN(n45) );
  AOI22_X1 U46 ( .A1(x[27]), .A2(net82897), .B1(y[27]), .B2(net83766), .ZN(n46) );
  AOI22_X1 U47 ( .A1(x[26]), .A2(net82897), .B1(y[26]), .B2(net83766), .ZN(n47) );
  AOI22_X1 U48 ( .A1(x[25]), .A2(net82897), .B1(y[25]), .B2(net94624), .ZN(n48) );
  AOI22_X1 U49 ( .A1(x[24]), .A2(net82897), .B1(y[24]), .B2(net83766), .ZN(n49) );
  AOI22_X1 U50 ( .A1(x[23]), .A2(net82897), .B1(y[23]), .B2(net83766), .ZN(n50) );
  AOI22_X1 U51 ( .A1(x[22]), .A2(net82897), .B1(y[22]), .B2(net83766), .ZN(n51) );
  AOI22_X1 U52 ( .A1(x[21]), .A2(net82897), .B1(y[21]), .B2(net83766), .ZN(n52) );
  AOI22_X1 U53 ( .A1(x[20]), .A2(net82897), .B1(y[20]), .B2(net83766), .ZN(n53) );
  AOI22_X1 U54 ( .A1(x[1]), .A2(net88219), .B1(net94624), .B2(y[1]), .ZN(n54)
         );
  AOI22_X1 U55 ( .A1(x[19]), .A2(net82897), .B1(y[19]), .B2(net83766), .ZN(n55) );
  AOI22_X1 U56 ( .A1(x[18]), .A2(net82897), .B1(y[18]), .B2(net83766), .ZN(n56) );
  AOI22_X1 U57 ( .A1(x[17]), .A2(net82897), .B1(y[17]), .B2(net83766), .ZN(n57) );
  AOI22_X1 U58 ( .A1(x[16]), .A2(net82897), .B1(y[16]), .B2(net83766), .ZN(n58) );
  AOI22_X1 U59 ( .A1(x[15]), .A2(net82700), .B1(net83357), .B2(y[15]), .ZN(n59) );
  AOI22_X1 U61 ( .A1(x[13]), .A2(net82700), .B1(net107657), .B2(y[13]), .ZN(
        n61) );
  AOI22_X1 U60 ( .A1(net76465), .A2(x[14]), .B1(y[14]), .B2(net83357), .ZN(n60) );
  AOI22_X1 U40 ( .A1(x[3]), .A2(net88219), .B1(y[3]), .B2(net75025), .ZN(n40)
         );
  AOI22_X1 U39 ( .A1(x[4]), .A2(net82700), .B1(y[4]), .B2(net107657), .ZN(n39)
         );
  AOI22_X1 U64 ( .A1(net75011), .A2(x[10]), .B1(net75023), .B2(y[10]), .ZN(n64) );
  AOI22_X1 U62 ( .A1(net112175), .A2(x[12]), .B1(net75023), .B2(y[12]), .ZN(
        n62) );
  AOI22_X1 U63 ( .A1(net75011), .A2(x[11]), .B1(net75023), .B2(y[11]), .ZN(n63) );
  AOI22_X1 U65 ( .A1(net76465), .A2(x[0]), .B1(net75015), .B2(y[0]), .ZN(n65)
         );
  AOI22_X1 U36 ( .A1(net112175), .A2(x[7]), .B1(net75015), .B2(y[7]), .ZN(n36)
         );
  AOI22_X1 U34 ( .A1(x[9]), .A2(net76465), .B1(net75015), .B2(y[9]), .ZN(n34)
         );
  INV_X1 U1 ( .A(n34), .ZN(net74051) );
  INV_X1 U5 ( .A(net75025), .ZN(net112175) );
  INV_X1 U8 ( .A(sel), .ZN(net75011) );
  INV_X1 U12 ( .A(n63), .ZN(net74053) );
  INV_X1 U14 ( .A(n62), .ZN(net74054) );
  CLKBUF_X1 U15 ( .A(net75011), .Z(net88219) );
  INV_X1 U16 ( .A(n37), .ZN(m[6]) );
  CLKBUF_X1 U17 ( .A(net75025), .Z(net94624) );
  INV_X1 U19 ( .A(n65), .ZN(net74042) );
  CLKBUF_X1 U20 ( .A(net94624), .Z(net83766) );
  INV_X1 U22 ( .A(net83766), .ZN(net82897) );
  INV_X1 U23 ( .A(n61), .ZN(m[13]) );
  INV_X1 U24 ( .A(n64), .ZN(net74052) );
  INV_X1 U25 ( .A(n35), .ZN(m[8]) );
  INV_X1 U26 ( .A(n60), .ZN(net74056) );
  INV_X1 U27 ( .A(n36), .ZN(net74049) );
  INV_X1 U28 ( .A(n38), .ZN(m[5]) );
  INV_X1 U29 ( .A(n54), .ZN(m[1]) );
  INV_X1 U30 ( .A(n40), .ZN(net74045) );
  INV_X1 U31 ( .A(n39), .ZN(net74046) );
  INV_X1 U32 ( .A(n58), .ZN(m[16]) );
  INV_X1 U33 ( .A(n52), .ZN(m[21]) );
  INV_X1 U66 ( .A(n53), .ZN(m[20]) );
  INV_X1 U67 ( .A(n55), .ZN(m[19]) );
  INV_X1 U68 ( .A(n57), .ZN(m[17]) );
  INV_X1 U69 ( .A(n56), .ZN(m[18]) );
  INV_X1 U70 ( .A(n42), .ZN(m[30]) );
  INV_X1 U71 ( .A(n45), .ZN(m[28]) );
  INV_X1 U72 ( .A(n46), .ZN(m[27]) );
  INV_X1 U73 ( .A(n48), .ZN(m[25]) );
  INV_X1 U74 ( .A(n47), .ZN(m[26]) );
  INV_X1 U75 ( .A(n41), .ZN(m[31]) );
  INV_X1 U76 ( .A(n51), .ZN(m[22]) );
  INV_X1 U77 ( .A(n50), .ZN(m[23]) );
  INV_X1 U78 ( .A(n44), .ZN(m[29]) );
  INV_X1 U79 ( .A(n49), .ZN(m[24]) );
  INV_X1 U80 ( .A(n59), .ZN(m[15]) );
  CLKBUF_X1 U2 ( .A(net75025), .Z(net75015) );
  BUF_X1 U3 ( .A(net75023), .Z(net107657) );
  CLKBUF_X1 U4 ( .A(net75011), .Z(net76465) );
  BUF_X1 U6 ( .A(net75011), .Z(net82700) );
  CLKBUF_X1 U7 ( .A(sel), .Z(net75025) );
  BUF_X2 U9 ( .A(sel), .Z(net75023) );
  INV_X1 U10 ( .A(n43), .ZN(m[2]) );
  BUF_X1 U11 ( .A(net75023), .Z(net83357) );
endmodule


module ALU_N32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n202, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78,
         n79, n81, n82, n84, n85, n86, n87, n88, n89, n91, n92, n94, n95, n96,
         n97, n98, n99, n101, n102, n104, n105, n106, n107, n108, n109, n111,
         n112, n114, n115, n116, n117, n118, n119, n121, n122, n124, n125,
         n126, n127, n128, n129, n131, n132, n134, n135, n136, n137, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n201, n93, n90, n83, n80, n73, n200,
         n138, n133, n130, n123, n120, n113, n110, n103, n100, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266;

  AOI21_X1 U65 ( .B1(n65), .B2(n204), .A(n66), .ZN(LE) );
  AOI22_X1 U66 ( .A1(A[30]), .A2(n237), .B1(n68), .B2(n69), .ZN(n67) );
  AOI21_X1 U67 ( .B1(n70), .B2(n71), .A(n72), .ZN(n68) );
  NAND2_X1 U69 ( .A1(n77), .A2(n78), .ZN(n74) );
  NAND2_X1 U72 ( .A1(n87), .A2(n88), .ZN(n84) );
  NAND2_X1 U75 ( .A1(n97), .A2(n98), .ZN(n94) );
  NAND2_X1 U78 ( .A1(n107), .A2(n108), .ZN(n104) );
  NAND2_X1 U81 ( .A1(n117), .A2(n118), .ZN(n114) );
  NAND2_X1 U84 ( .A1(n127), .A2(n128), .ZN(n124) );
  OAI21_X1 U89 ( .B1(n234), .B2(n141), .A(B[1]), .ZN(n139) );
  NAND2_X1 U90 ( .A1(A[0]), .A2(n266), .ZN(n141) );
  NOR2_X1 U91 ( .A1(n142), .A2(n143), .ZN(n129) );
  NOR2_X1 U92 ( .A1(n144), .A2(n145), .ZN(n119) );
  NOR2_X1 U93 ( .A1(n146), .A2(n147), .ZN(n109) );
  NOR2_X1 U94 ( .A1(n148), .A2(n149), .ZN(n99) );
  NOR2_X1 U95 ( .A1(n150), .A2(n151), .ZN(n89) );
  NOR2_X1 U96 ( .A1(n152), .A2(n153), .ZN(n79) );
  NOR2_X1 U97 ( .A1(n154), .A2(n155), .ZN(n70) );
  OAI21_X1 U98 ( .B1(n66), .B2(n156), .A(n65), .ZN(n202) );
  NAND2_X1 U99 ( .A1(A[31]), .A2(n236), .ZN(n65) );
  AOI22_X1 U100 ( .A1(B[30]), .A2(n205), .B1(n157), .B2(n69), .ZN(n156) );
  XOR2_X1 U101 ( .A(n205), .B(B[30]), .Z(n69) );
  AOI21_X1 U102 ( .B1(n158), .B2(n206), .A(n155), .ZN(n157) );
  NOR2_X1 U104 ( .A1(n238), .A2(A[29]), .ZN(n72) );
  AOI21_X1 U105 ( .B1(n159), .B2(n76), .A(n160), .ZN(n158) );
  NOR2_X1 U106 ( .A1(n160), .A2(n154), .ZN(n76) );
  NOR2_X1 U108 ( .A1(n239), .A2(A[28]), .ZN(n160) );
  AOI21_X1 U109 ( .B1(n161), .B2(n75), .A(n207), .ZN(n159) );
  NAND2_X1 U110 ( .A1(A[27]), .A2(n240), .ZN(n77) );
  OR2_X1 U111 ( .A1(n240), .A2(A[27]), .ZN(n75) );
  AOI21_X1 U112 ( .B1(n162), .B2(n208), .A(n163), .ZN(n161) );
  NAND2_X1 U113 ( .A1(n209), .A2(n78), .ZN(n81) );
  NAND2_X1 U114 ( .A1(A[26]), .A2(n241), .ZN(n78) );
  NOR2_X1 U115 ( .A1(n241), .A2(A[26]), .ZN(n163) );
  AOI21_X1 U116 ( .B1(n164), .B2(n210), .A(n153), .ZN(n162) );
  NOR2_X1 U118 ( .A1(n242), .A2(A[25]), .ZN(n82) );
  AOI21_X1 U119 ( .B1(n165), .B2(n86), .A(n166), .ZN(n164) );
  NOR2_X1 U120 ( .A1(n166), .A2(n152), .ZN(n86) );
  NOR2_X1 U122 ( .A1(n243), .A2(A[24]), .ZN(n166) );
  AOI21_X1 U123 ( .B1(n167), .B2(n85), .A(n211), .ZN(n165) );
  NAND2_X1 U124 ( .A1(A[23]), .A2(n244), .ZN(n87) );
  OR2_X1 U125 ( .A1(n244), .A2(A[23]), .ZN(n85) );
  AOI21_X1 U126 ( .B1(n168), .B2(n212), .A(n169), .ZN(n167) );
  NAND2_X1 U127 ( .A1(n213), .A2(n88), .ZN(n91) );
  NAND2_X1 U128 ( .A1(A[22]), .A2(n245), .ZN(n88) );
  NOR2_X1 U129 ( .A1(n245), .A2(A[22]), .ZN(n169) );
  AOI21_X1 U130 ( .B1(n170), .B2(n214), .A(n151), .ZN(n168) );
  NOR2_X1 U132 ( .A1(n246), .A2(A[21]), .ZN(n92) );
  AOI21_X1 U133 ( .B1(n171), .B2(n96), .A(n172), .ZN(n170) );
  NOR2_X1 U134 ( .A1(n172), .A2(n150), .ZN(n96) );
  NOR2_X1 U136 ( .A1(n247), .A2(A[20]), .ZN(n172) );
  AOI21_X1 U137 ( .B1(n173), .B2(n95), .A(n215), .ZN(n171) );
  NAND2_X1 U138 ( .A1(A[19]), .A2(n248), .ZN(n97) );
  OR2_X1 U139 ( .A1(n248), .A2(A[19]), .ZN(n95) );
  AOI21_X1 U140 ( .B1(n174), .B2(n216), .A(n175), .ZN(n173) );
  NAND2_X1 U141 ( .A1(n217), .A2(n98), .ZN(n101) );
  NAND2_X1 U142 ( .A1(A[18]), .A2(n249), .ZN(n98) );
  NOR2_X1 U143 ( .A1(n249), .A2(A[18]), .ZN(n175) );
  AOI21_X1 U144 ( .B1(n176), .B2(n218), .A(n149), .ZN(n174) );
  NOR2_X1 U146 ( .A1(n250), .A2(A[17]), .ZN(n102) );
  AOI21_X1 U147 ( .B1(n177), .B2(n106), .A(n178), .ZN(n176) );
  NOR2_X1 U148 ( .A1(n178), .A2(n148), .ZN(n106) );
  NOR2_X1 U150 ( .A1(n251), .A2(A[16]), .ZN(n178) );
  AOI21_X1 U151 ( .B1(n179), .B2(n105), .A(n219), .ZN(n177) );
  NAND2_X1 U152 ( .A1(A[15]), .A2(n252), .ZN(n107) );
  OR2_X1 U153 ( .A1(n252), .A2(A[15]), .ZN(n105) );
  AOI21_X1 U154 ( .B1(n180), .B2(n220), .A(n181), .ZN(n179) );
  NAND2_X1 U155 ( .A1(n221), .A2(n108), .ZN(n111) );
  NAND2_X1 U156 ( .A1(A[14]), .A2(n253), .ZN(n108) );
  NOR2_X1 U157 ( .A1(n253), .A2(A[14]), .ZN(n181) );
  AOI21_X1 U158 ( .B1(n182), .B2(n222), .A(n147), .ZN(n180) );
  NOR2_X1 U160 ( .A1(n254), .A2(A[13]), .ZN(n112) );
  AOI21_X1 U161 ( .B1(n183), .B2(n116), .A(n184), .ZN(n182) );
  NOR2_X1 U162 ( .A1(n184), .A2(n146), .ZN(n116) );
  NOR2_X1 U164 ( .A1(n255), .A2(A[12]), .ZN(n184) );
  AOI21_X1 U165 ( .B1(n185), .B2(n115), .A(n223), .ZN(n183) );
  NAND2_X1 U166 ( .A1(A[11]), .A2(n256), .ZN(n117) );
  OR2_X1 U167 ( .A1(n256), .A2(A[11]), .ZN(n115) );
  AOI21_X1 U168 ( .B1(n186), .B2(n224), .A(n187), .ZN(n185) );
  NAND2_X1 U169 ( .A1(n225), .A2(n118), .ZN(n121) );
  NAND2_X1 U170 ( .A1(A[10]), .A2(n257), .ZN(n118) );
  NOR2_X1 U171 ( .A1(n257), .A2(A[10]), .ZN(n187) );
  AOI21_X1 U172 ( .B1(n188), .B2(n226), .A(n145), .ZN(n186) );
  NOR2_X1 U174 ( .A1(n258), .A2(A[9]), .ZN(n122) );
  AOI21_X1 U175 ( .B1(n189), .B2(n126), .A(n190), .ZN(n188) );
  NOR2_X1 U176 ( .A1(n190), .A2(n144), .ZN(n126) );
  NOR2_X1 U178 ( .A1(n259), .A2(A[8]), .ZN(n190) );
  AOI21_X1 U179 ( .B1(n191), .B2(n125), .A(n227), .ZN(n189) );
  NAND2_X1 U180 ( .A1(A[7]), .A2(n260), .ZN(n127) );
  OR2_X1 U181 ( .A1(n260), .A2(A[7]), .ZN(n125) );
  AOI21_X1 U182 ( .B1(n192), .B2(n228), .A(n193), .ZN(n191) );
  NAND2_X1 U183 ( .A1(n229), .A2(n128), .ZN(n131) );
  NAND2_X1 U184 ( .A1(A[6]), .A2(n261), .ZN(n128) );
  NOR2_X1 U185 ( .A1(n261), .A2(A[6]), .ZN(n193) );
  AOI21_X1 U186 ( .B1(n194), .B2(n230), .A(n143), .ZN(n192) );
  NOR2_X1 U188 ( .A1(n262), .A2(A[5]), .ZN(n132) );
  AOI21_X1 U189 ( .B1(n195), .B2(n135), .A(n196), .ZN(n194) );
  NOR2_X1 U190 ( .A1(n196), .A2(n142), .ZN(n135) );
  NOR2_X1 U192 ( .A1(n263), .A2(A[4]), .ZN(n196) );
  AOI21_X1 U193 ( .B1(n197), .B2(n134), .A(n231), .ZN(n195) );
  NAND2_X1 U194 ( .A1(A[3]), .A2(n264), .ZN(n136) );
  OR2_X1 U195 ( .A1(n264), .A2(A[3]), .ZN(n134) );
  AOI21_X1 U196 ( .B1(n233), .B2(n140), .A(n198), .ZN(n197) );
  NOR2_X1 U197 ( .A1(n198), .A2(n232), .ZN(n140) );
  NAND2_X1 U198 ( .A1(A[2]), .A2(n265), .ZN(n137) );
  NOR2_X1 U199 ( .A1(n265), .A2(A[2]), .ZN(n198) );
  NOR2_X1 U202 ( .A1(n266), .A2(A[0]), .ZN(n201) );
  NOR2_X1 U203 ( .A1(n236), .A2(A[31]), .ZN(n66) );
  INV_X1 U1 ( .A(n121), .ZN(n224) );
  INV_X1 U2 ( .A(n101), .ZN(n216) );
  INV_X1 U3 ( .A(n81), .ZN(n208) );
  INV_X1 U4 ( .A(n137), .ZN(n232) );
  INV_X1 U5 ( .A(n111), .ZN(n220) );
  INV_X1 U6 ( .A(n112), .ZN(n222) );
  INV_X1 U7 ( .A(n91), .ZN(n212) );
  INV_X1 U8 ( .A(n92), .ZN(n214) );
  INV_X1 U9 ( .A(n117), .ZN(n223) );
  INV_X1 U10 ( .A(n97), .ZN(n215) );
  INV_X1 U11 ( .A(n131), .ZN(n228) );
  INV_X1 U12 ( .A(n132), .ZN(n230) );
  INV_X1 U13 ( .A(n122), .ZN(n226) );
  INV_X1 U14 ( .A(n102), .ZN(n218) );
  INV_X1 U15 ( .A(n82), .ZN(n210) );
  INV_X1 U16 ( .A(n77), .ZN(n207) );
  INV_X1 U17 ( .A(n193), .ZN(n229) );
  INV_X1 U18 ( .A(n187), .ZN(n225) );
  INV_X1 U19 ( .A(n181), .ZN(n221) );
  INV_X1 U20 ( .A(n127), .ZN(n227) );
  INV_X1 U21 ( .A(n175), .ZN(n217) );
  INV_X1 U22 ( .A(n169), .ZN(n213) );
  INV_X1 U23 ( .A(n163), .ZN(n209) );
  INV_X1 U24 ( .A(n72), .ZN(n206) );
  INV_X1 U25 ( .A(n107), .ZN(n219) );
  INV_X1 U26 ( .A(n87), .ZN(n211) );
  INV_X1 U27 ( .A(n136), .ZN(n231) );
  INV_X1 U28 ( .A(B[4]), .ZN(n263) );
  INV_X1 U29 ( .A(n67), .ZN(n204) );
  INV_X1 U30 ( .A(B[0]), .ZN(n266) );
  INV_X1 U31 ( .A(B[3]), .ZN(n264) );
  INV_X1 U32 ( .A(B[15]), .ZN(n252) );
  INV_X1 U33 ( .A(A[30]), .ZN(n205) );
  INV_X1 U34 ( .A(n141), .ZN(n235) );
  INV_X1 U35 ( .A(A[1]), .ZN(n234) );
  INV_X1 U36 ( .A(B[2]), .ZN(n265) );
  INV_X1 U37 ( .A(B[9]), .ZN(n258) );
  INV_X1 U38 ( .A(B[12]), .ZN(n255) );
  INV_X1 U39 ( .A(B[14]), .ZN(n253) );
  INV_X1 U40 ( .A(B[8]), .ZN(n259) );
  INV_X1 U41 ( .A(B[5]), .ZN(n262) );
  INV_X1 U42 ( .A(B[6]), .ZN(n261) );
  INV_X1 U43 ( .A(B[10]), .ZN(n257) );
  INV_X1 U44 ( .A(B[11]), .ZN(n256) );
  INV_X1 U45 ( .A(B[7]), .ZN(n260) );
  INV_X1 U46 ( .A(n202), .ZN(GE) );
  INV_X1 U47 ( .A(n199), .ZN(n233) );
  INV_X1 U48 ( .A(B[13]), .ZN(n254) );
  INV_X1 U49 ( .A(B[28]), .ZN(n239) );
  INV_X1 U50 ( .A(B[25]), .ZN(n242) );
  INV_X1 U51 ( .A(B[26]), .ZN(n241) );
  INV_X1 U52 ( .A(B[31]), .ZN(n236) );
  INV_X1 U53 ( .A(B[21]), .ZN(n246) );
  INV_X1 U54 ( .A(B[20]), .ZN(n247) );
  INV_X1 U55 ( .A(B[17]), .ZN(n250) );
  INV_X1 U56 ( .A(B[16]), .ZN(n251) );
  INV_X1 U57 ( .A(B[18]), .ZN(n249) );
  INV_X1 U58 ( .A(B[29]), .ZN(n238) );
  INV_X1 U59 ( .A(B[22]), .ZN(n245) );
  INV_X1 U60 ( .A(B[24]), .ZN(n243) );
  INV_X1 U61 ( .A(B[27]), .ZN(n240) );
  INV_X1 U62 ( .A(B[19]), .ZN(n248) );
  INV_X1 U63 ( .A(B[23]), .ZN(n244) );
  INV_X1 U64 ( .A(B[30]), .ZN(n237) );
  AND2_X1 U68 ( .A1(A[4]), .A2(n263), .ZN(n142) );
  AND2_X1 U70 ( .A1(A[5]), .A2(n262), .ZN(n143) );
  OAI211_X1 U71 ( .C1(A[1]), .C2(n235), .A(n139), .B(n140), .ZN(n138) );
  AND2_X1 U73 ( .A1(A[13]), .A2(n254), .ZN(n147) );
  AND2_X1 U74 ( .A1(A[12]), .A2(n255), .ZN(n146) );
  AOI211_X1 U76 ( .C1(n119), .C2(n120), .A(n121), .B(n122), .ZN(n113) );
  OAI211_X1 U77 ( .C1(n123), .C2(n124), .A(n125), .B(n126), .ZN(n120) );
  AND2_X1 U79 ( .A1(A[21]), .A2(n246), .ZN(n151) );
  AND2_X1 U80 ( .A1(A[20]), .A2(n247), .ZN(n150) );
  AOI211_X1 U82 ( .C1(n99), .C2(n100), .A(n101), .B(n102), .ZN(n93) );
  OAI211_X1 U83 ( .C1(n103), .C2(n104), .A(n105), .B(n106), .ZN(n100) );
  AOI211_X1 U85 ( .C1(n79), .C2(n80), .A(n81), .B(n82), .ZN(n73) );
  OAI211_X1 U86 ( .C1(n83), .C2(n84), .A(n85), .B(n86), .ZN(n80) );
  OAI22_X1 U87 ( .A1(n200), .A2(B[1]), .B1(n234), .B2(n201), .ZN(n199) );
  AND2_X1 U88 ( .A1(n201), .A2(n234), .ZN(n200) );
  AND2_X1 U103 ( .A1(A[8]), .A2(n259), .ZN(n144) );
  AND2_X1 U107 ( .A1(A[9]), .A2(n258), .ZN(n145) );
  AOI211_X1 U117 ( .C1(n129), .C2(n130), .A(n131), .B(n132), .ZN(n123) );
  NAND3_X1 U121 ( .A1(n133), .A2(n134), .A3(n135), .ZN(n130) );
  NAND3_X1 U131 ( .A1(n136), .A2(n137), .A3(n138), .ZN(n133) );
  AND2_X1 U135 ( .A1(A[17]), .A2(n250), .ZN(n149) );
  AND2_X1 U145 ( .A1(A[16]), .A2(n251), .ZN(n148) );
  AOI211_X1 U149 ( .C1(n109), .C2(n110), .A(n111), .B(n112), .ZN(n103) );
  OAI211_X1 U159 ( .C1(n113), .C2(n114), .A(n115), .B(n116), .ZN(n110) );
  AND2_X1 U163 ( .A1(A[24]), .A2(n243), .ZN(n152) );
  AND2_X1 U173 ( .A1(A[25]), .A2(n242), .ZN(n153) );
  AOI211_X1 U177 ( .C1(n89), .C2(n90), .A(n91), .B(n92), .ZN(n83) );
  OAI211_X1 U187 ( .C1(n93), .C2(n94), .A(n95), .B(n96), .ZN(n90) );
  AND2_X1 U191 ( .A1(A[28]), .A2(n239), .ZN(n154) );
  AND2_X1 U200 ( .A1(A[29]), .A2(n238), .ZN(n155) );
  OAI211_X1 U201 ( .C1(n73), .C2(n74), .A(n75), .B(n76), .ZN(n71) );
endmodule


module ALU_N32_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n202, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n161, n162, n163, n164, n167, n168, n169, n170, n173, n174, n175,
         n176, n179, n180, n181, n182, n185, n186, n187, n188, n191, n192,
         n193, n194, n197, n198, n200, n201, n199, n196, n195, n190, n189,
         n184, n183, n178, n177, n172, n171, n166, n165, n160, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265;

  AOI21_X1 U65 ( .B1(n65), .B2(n204), .A(n66), .ZN(GE) );
  AOI22_X1 U66 ( .A1(B[30]), .A2(n205), .B1(n68), .B2(n69), .ZN(n67) );
  AOI21_X1 U67 ( .B1(n70), .B2(n71), .A(n72), .ZN(n68) );
  AOI21_X1 U68 ( .B1(n73), .B2(n74), .A(n75), .ZN(n70) );
  AOI21_X1 U69 ( .B1(n76), .B2(n77), .A(n78), .ZN(n73) );
  AOI21_X1 U70 ( .B1(n79), .B2(n212), .A(n211), .ZN(n76) );
  AOI21_X1 U71 ( .B1(n82), .B2(n83), .A(n84), .ZN(n79) );
  AOI21_X1 U72 ( .B1(n85), .B2(n86), .A(n87), .ZN(n82) );
  AOI21_X1 U73 ( .B1(n88), .B2(n89), .A(n90), .ZN(n85) );
  AOI21_X1 U74 ( .B1(n91), .B2(n220), .A(n219), .ZN(n88) );
  AOI21_X1 U75 ( .B1(n94), .B2(n95), .A(n96), .ZN(n91) );
  AOI21_X1 U76 ( .B1(n97), .B2(n98), .A(n99), .ZN(n94) );
  AOI21_X1 U77 ( .B1(n100), .B2(n101), .A(n102), .ZN(n97) );
  AOI21_X1 U78 ( .B1(n103), .B2(n228), .A(n227), .ZN(n100) );
  AOI21_X1 U79 ( .B1(n106), .B2(n107), .A(n108), .ZN(n103) );
  AOI21_X1 U80 ( .B1(n109), .B2(n110), .A(n111), .ZN(n106) );
  AOI21_X1 U81 ( .B1(n112), .B2(n113), .A(n114), .ZN(n109) );
  AOI21_X1 U82 ( .B1(n115), .B2(n236), .A(n235), .ZN(n112) );
  AOI21_X1 U83 ( .B1(n118), .B2(n119), .A(n120), .ZN(n115) );
  AOI21_X1 U84 ( .B1(n121), .B2(n122), .A(n123), .ZN(n118) );
  AOI21_X1 U85 ( .B1(n124), .B2(n125), .A(n126), .ZN(n121) );
  AOI21_X1 U86 ( .B1(n127), .B2(n244), .A(n243), .ZN(n124) );
  AOI21_X1 U87 ( .B1(n130), .B2(n131), .A(n132), .ZN(n127) );
  AOI21_X1 U88 ( .B1(n133), .B2(n134), .A(n135), .ZN(n130) );
  AOI21_X1 U89 ( .B1(n136), .B2(n137), .A(n138), .ZN(n133) );
  AOI21_X1 U90 ( .B1(n139), .B2(n252), .A(n251), .ZN(n136) );
  AOI21_X1 U91 ( .B1(n142), .B2(n143), .A(n144), .ZN(n139) );
  AOI21_X1 U92 ( .B1(n145), .B2(n146), .A(n147), .ZN(n142) );
  AOI21_X1 U93 ( .B1(n148), .B2(n149), .A(n150), .ZN(n145) );
  AOI21_X1 U94 ( .B1(n151), .B2(n152), .A(n259), .ZN(n148) );
  AOI22_X1 U95 ( .A1(n154), .A2(n265), .B1(A[1]), .B2(n155), .ZN(n151) );
  OR2_X1 U96 ( .A1(n155), .A2(A[1]), .ZN(n154) );
  NAND2_X1 U97 ( .A1(B[0]), .A2(n262), .ZN(n155) );
  OAI21_X1 U98 ( .B1(n66), .B2(n156), .A(n65), .ZN(n202) );
  NAND2_X1 U99 ( .A1(A[31]), .A2(n263), .ZN(n65) );
  AOI22_X1 U100 ( .A1(A[30]), .A2(n264), .B1(n157), .B2(n69), .ZN(n156) );
  XOR2_X1 U101 ( .A(A[30]), .B(n264), .Z(n69) );
  AOI21_X1 U102 ( .B1(n158), .B2(n159), .A(n206), .ZN(n157) );
  NAND2_X1 U103 ( .A1(B[29]), .A2(n207), .ZN(n71) );
  NOR2_X1 U105 ( .A1(n162), .A2(n75), .ZN(n74) );
  NAND2_X1 U107 ( .A1(B[27]), .A2(n210), .ZN(n77) );
  NAND2_X1 U108 ( .A1(n209), .A2(n163), .ZN(n161) );
  NOR2_X1 U109 ( .A1(n210), .A2(B[27]), .ZN(n78) );
  NAND2_X1 U111 ( .A1(B[25]), .A2(n215), .ZN(n83) );
  NAND2_X1 U112 ( .A1(n163), .A2(n80), .ZN(n81) );
  NAND2_X1 U113 ( .A1(B[26]), .A2(n213), .ZN(n80) );
  OR2_X1 U114 ( .A1(n213), .A2(B[26]), .ZN(n163) );
  NOR2_X1 U116 ( .A1(n168), .A2(n87), .ZN(n86) );
  NAND2_X1 U118 ( .A1(B[23]), .A2(n218), .ZN(n89) );
  NAND2_X1 U119 ( .A1(n217), .A2(n169), .ZN(n167) );
  NOR2_X1 U120 ( .A1(n218), .A2(B[23]), .ZN(n90) );
  NAND2_X1 U122 ( .A1(B[21]), .A2(n223), .ZN(n95) );
  NAND2_X1 U123 ( .A1(n169), .A2(n92), .ZN(n93) );
  NAND2_X1 U124 ( .A1(B[22]), .A2(n221), .ZN(n92) );
  OR2_X1 U125 ( .A1(n221), .A2(B[22]), .ZN(n169) );
  NOR2_X1 U127 ( .A1(n174), .A2(n99), .ZN(n98) );
  NAND2_X1 U129 ( .A1(B[19]), .A2(n226), .ZN(n101) );
  NAND2_X1 U130 ( .A1(n225), .A2(n175), .ZN(n173) );
  NOR2_X1 U131 ( .A1(n226), .A2(B[19]), .ZN(n102) );
  NAND2_X1 U133 ( .A1(B[17]), .A2(n231), .ZN(n107) );
  NAND2_X1 U134 ( .A1(n175), .A2(n104), .ZN(n105) );
  NAND2_X1 U135 ( .A1(B[18]), .A2(n229), .ZN(n104) );
  OR2_X1 U136 ( .A1(n229), .A2(B[18]), .ZN(n175) );
  NOR2_X1 U138 ( .A1(n180), .A2(n111), .ZN(n110) );
  NAND2_X1 U140 ( .A1(B[15]), .A2(n234), .ZN(n113) );
  NAND2_X1 U141 ( .A1(n233), .A2(n181), .ZN(n179) );
  NOR2_X1 U142 ( .A1(n234), .A2(B[15]), .ZN(n114) );
  NAND2_X1 U144 ( .A1(B[13]), .A2(n239), .ZN(n119) );
  NAND2_X1 U145 ( .A1(n181), .A2(n116), .ZN(n117) );
  NAND2_X1 U146 ( .A1(B[14]), .A2(n237), .ZN(n116) );
  OR2_X1 U147 ( .A1(n237), .A2(B[14]), .ZN(n181) );
  NOR2_X1 U149 ( .A1(n186), .A2(n123), .ZN(n122) );
  NAND2_X1 U151 ( .A1(B[11]), .A2(n242), .ZN(n125) );
  NAND2_X1 U152 ( .A1(n241), .A2(n187), .ZN(n185) );
  NOR2_X1 U153 ( .A1(n242), .A2(B[11]), .ZN(n126) );
  NAND2_X1 U155 ( .A1(B[9]), .A2(n247), .ZN(n131) );
  NAND2_X1 U156 ( .A1(n187), .A2(n128), .ZN(n129) );
  NAND2_X1 U157 ( .A1(B[10]), .A2(n245), .ZN(n128) );
  OR2_X1 U158 ( .A1(n245), .A2(B[10]), .ZN(n187) );
  NOR2_X1 U160 ( .A1(n192), .A2(n135), .ZN(n134) );
  NAND2_X1 U162 ( .A1(B[7]), .A2(n250), .ZN(n137) );
  NAND2_X1 U163 ( .A1(n249), .A2(n193), .ZN(n191) );
  NOR2_X1 U164 ( .A1(n250), .A2(B[7]), .ZN(n138) );
  NAND2_X1 U166 ( .A1(B[5]), .A2(n255), .ZN(n143) );
  NAND2_X1 U167 ( .A1(n193), .A2(n140), .ZN(n141) );
  NAND2_X1 U168 ( .A1(B[6]), .A2(n253), .ZN(n140) );
  OR2_X1 U169 ( .A1(n253), .A2(B[6]), .ZN(n193) );
  NOR2_X1 U171 ( .A1(n197), .A2(n147), .ZN(n146) );
  NAND2_X1 U173 ( .A1(B[3]), .A2(n258), .ZN(n149) );
  NAND2_X1 U177 ( .A1(B[2]), .A2(n260), .ZN(n153) );
  AOI21_X1 U178 ( .B1(A[1]), .B2(n200), .A(n265), .ZN(n201) );
  NOR2_X1 U179 ( .A1(n262), .A2(B[0]), .ZN(n200) );
  OR2_X1 U180 ( .A1(n260), .A2(B[2]), .ZN(n198) );
  NOR2_X1 U181 ( .A1(n258), .A2(B[3]), .ZN(n150) );
  NOR2_X1 U182 ( .A1(n197), .A2(n144), .ZN(n194) );
  NOR2_X1 U183 ( .A1(n255), .A2(B[5]), .ZN(n144) );
  NOR2_X1 U184 ( .A1(n256), .A2(B[4]), .ZN(n197) );
  NOR2_X1 U185 ( .A1(n192), .A2(n132), .ZN(n188) );
  NOR2_X1 U186 ( .A1(n247), .A2(B[9]), .ZN(n132) );
  NOR2_X1 U187 ( .A1(n248), .A2(B[8]), .ZN(n192) );
  NOR2_X1 U188 ( .A1(n186), .A2(n120), .ZN(n182) );
  NOR2_X1 U189 ( .A1(n239), .A2(B[13]), .ZN(n120) );
  NOR2_X1 U190 ( .A1(n240), .A2(B[12]), .ZN(n186) );
  NOR2_X1 U191 ( .A1(n180), .A2(n108), .ZN(n176) );
  NOR2_X1 U192 ( .A1(n231), .A2(B[17]), .ZN(n108) );
  NOR2_X1 U193 ( .A1(n232), .A2(B[16]), .ZN(n180) );
  NOR2_X1 U194 ( .A1(n174), .A2(n96), .ZN(n170) );
  NOR2_X1 U195 ( .A1(n223), .A2(B[21]), .ZN(n96) );
  NOR2_X1 U196 ( .A1(n224), .A2(B[20]), .ZN(n174) );
  NOR2_X1 U197 ( .A1(n168), .A2(n84), .ZN(n164) );
  NOR2_X1 U198 ( .A1(n215), .A2(B[25]), .ZN(n84) );
  NOR2_X1 U199 ( .A1(n216), .A2(B[24]), .ZN(n168) );
  NOR2_X1 U200 ( .A1(n162), .A2(n72), .ZN(n158) );
  NOR2_X1 U201 ( .A1(n207), .A2(B[29]), .ZN(n72) );
  NOR2_X1 U202 ( .A1(n208), .A2(B[28]), .ZN(n162) );
  NOR2_X1 U203 ( .A1(n263), .A2(A[31]), .ZN(n66) );
  INV_X1 U2 ( .A(n141), .ZN(n252) );
  INV_X1 U3 ( .A(n129), .ZN(n244) );
  INV_X1 U4 ( .A(n117), .ZN(n236) );
  INV_X1 U5 ( .A(n105), .ZN(n228) );
  INV_X1 U6 ( .A(n93), .ZN(n220) );
  INV_X1 U7 ( .A(n81), .ZN(n212) );
  INV_X1 U8 ( .A(n138), .ZN(n249) );
  INV_X1 U9 ( .A(n126), .ZN(n241) );
  INV_X1 U10 ( .A(n114), .ZN(n233) );
  INV_X1 U11 ( .A(n102), .ZN(n225) );
  INV_X1 U12 ( .A(n202), .ZN(LE) );
  INV_X1 U13 ( .A(A[0]), .ZN(n262) );
  INV_X1 U14 ( .A(A[7]), .ZN(n250) );
  INV_X1 U15 ( .A(A[11]), .ZN(n242) );
  INV_X1 U16 ( .A(A[8]), .ZN(n248) );
  INV_X1 U17 ( .A(A[9]), .ZN(n247) );
  INV_X1 U18 ( .A(A[5]), .ZN(n255) );
  INV_X1 U19 ( .A(n90), .ZN(n217) );
  INV_X1 U20 ( .A(n78), .ZN(n209) );
  INV_X1 U21 ( .A(A[12]), .ZN(n240) );
  INV_X1 U22 ( .A(A[3]), .ZN(n258) );
  INV_X1 U23 ( .A(A[4]), .ZN(n256) );
  INV_X1 U24 ( .A(A[6]), .ZN(n253) );
  INV_X1 U25 ( .A(A[10]), .ZN(n245) );
  INV_X1 U26 ( .A(A[2]), .ZN(n260) );
  INV_X1 U27 ( .A(n153), .ZN(n259) );
  INV_X1 U28 ( .A(n131), .ZN(n246) );
  INV_X1 U29 ( .A(n143), .ZN(n254) );
  INV_X1 U30 ( .A(n140), .ZN(n251) );
  INV_X1 U31 ( .A(A[15]), .ZN(n234) );
  INV_X1 U32 ( .A(A[16]), .ZN(n232) );
  INV_X1 U33 ( .A(A[28]), .ZN(n208) );
  INV_X1 U34 ( .A(A[17]), .ZN(n231) );
  INV_X1 U35 ( .A(A[21]), .ZN(n223) );
  INV_X1 U36 ( .A(A[25]), .ZN(n215) );
  INV_X1 U37 ( .A(A[27]), .ZN(n210) );
  INV_X1 U38 ( .A(A[20]), .ZN(n224) );
  INV_X1 U39 ( .A(A[24]), .ZN(n216) );
  INV_X1 U40 ( .A(A[13]), .ZN(n239) );
  INV_X1 U41 ( .A(A[29]), .ZN(n207) );
  INV_X1 U42 ( .A(A[19]), .ZN(n226) );
  INV_X1 U43 ( .A(A[23]), .ZN(n218) );
  INV_X1 U44 ( .A(A[18]), .ZN(n229) );
  INV_X1 U45 ( .A(A[22]), .ZN(n221) );
  INV_X1 U46 ( .A(A[26]), .ZN(n213) );
  INV_X1 U47 ( .A(A[14]), .ZN(n237) );
  INV_X1 U48 ( .A(n119), .ZN(n238) );
  INV_X1 U49 ( .A(n116), .ZN(n235) );
  INV_X1 U50 ( .A(n83), .ZN(n214) );
  INV_X1 U51 ( .A(n128), .ZN(n243) );
  INV_X1 U52 ( .A(n80), .ZN(n211) );
  INV_X1 U53 ( .A(n95), .ZN(n222) );
  INV_X1 U54 ( .A(n107), .ZN(n230) );
  INV_X1 U55 ( .A(n104), .ZN(n227) );
  INV_X1 U56 ( .A(n92), .ZN(n219) );
  INV_X1 U57 ( .A(n71), .ZN(n206) );
  INV_X1 U58 ( .A(n67), .ZN(n204) );
  INV_X1 U59 ( .A(A[30]), .ZN(n205) );
  INV_X1 U60 ( .A(n201), .ZN(n261) );
  INV_X1 U61 ( .A(n150), .ZN(n257) );
  INV_X1 U62 ( .A(B[1]), .ZN(n265) );
  INV_X1 U63 ( .A(B[30]), .ZN(n264) );
  INV_X1 U64 ( .A(B[31]), .ZN(n263) );
  OAI211_X1 U1 ( .C1(n190), .C2(n191), .A(n137), .B(n134), .ZN(n189) );
  AOI211_X1 U104 ( .C1(n194), .C2(n195), .A(n141), .B(n254), .ZN(n190) );
  OAI211_X1 U106 ( .C1(n178), .C2(n179), .A(n113), .B(n110), .ZN(n177) );
  AOI211_X1 U110 ( .C1(n182), .C2(n183), .A(n117), .B(n238), .ZN(n178) );
  OAI211_X1 U115 ( .C1(n166), .C2(n167), .A(n89), .B(n86), .ZN(n165) );
  AOI211_X1 U117 ( .C1(n170), .C2(n171), .A(n93), .B(n222), .ZN(n166) );
  NAND3_X1 U121 ( .A1(n196), .A2(n149), .A3(n146), .ZN(n195) );
  NAND3_X1 U126 ( .A1(n257), .A2(n198), .A3(n199), .ZN(n196) );
  OAI211_X1 U128 ( .C1(A[1]), .C2(n200), .A(n261), .B(n152), .ZN(n199) );
  AND2_X1 U132 ( .A1(B[4]), .A2(n256), .ZN(n147) );
  AND2_X1 U137 ( .A1(n198), .A2(n153), .ZN(n152) );
  AND2_X1 U139 ( .A1(B[8]), .A2(n248), .ZN(n135) );
  OAI211_X1 U143 ( .C1(n184), .C2(n185), .A(n125), .B(n122), .ZN(n183) );
  AOI211_X1 U148 ( .C1(n188), .C2(n189), .A(n129), .B(n246), .ZN(n184) );
  AND2_X1 U150 ( .A1(B[12]), .A2(n240), .ZN(n123) );
  AND2_X1 U154 ( .A1(B[16]), .A2(n232), .ZN(n111) );
  OAI211_X1 U159 ( .C1(n172), .C2(n173), .A(n101), .B(n98), .ZN(n171) );
  AOI211_X1 U161 ( .C1(n176), .C2(n177), .A(n105), .B(n230), .ZN(n172) );
  AND2_X1 U165 ( .A1(B[20]), .A2(n224), .ZN(n99) );
  AND2_X1 U170 ( .A1(B[24]), .A2(n216), .ZN(n87) );
  OAI211_X1 U172 ( .C1(n160), .C2(n161), .A(n77), .B(n74), .ZN(n159) );
  AOI211_X1 U174 ( .C1(n164), .C2(n165), .A(n81), .B(n214), .ZN(n160) );
  AND2_X1 U175 ( .A1(B[28]), .A2(n208), .ZN(n75) );
  AND2_X1 U176 ( .A1(LE), .A2(GE), .ZN(EQ) );
endmodule


module ALU_N32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] ,
         \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n97, n104, n111, n112,
         n114, n115, n118, n122, n125, n129, n136, n140, n141, net82621,
         net83063, net83123, net83718, net84366, net84352, net84350, net84349,
         net84344, net84329, net84304, net84303, net84298, net84293, net86108,
         net88213, net88223, net95093, net95224, net95222, net97351, net99106,
         net99092, net99109, net99128, net99126, net99137, net99158, net74518,
         net110243, net110231, net110228, net110223, net74529, n93, n91,
         net112065, net112146, net112161, net112169, net112166, net116127,
         net116123, net116117, net116113, net116111, net116094, net116079,
         net116070, net116138, net99183, net95223, net95128, net95052,
         net124940, net124943, net125026, net125034, net82778, n89, net112093,
         net112060, net112059, net112050, net110245, net95236, net95234,
         net95098, net99082, net99050, net97413, net95122, net95089, net125041,
         net125031, net116155, net116153, net84338, net110221, net110220,
         net110131, net99166, net125015, net125007, net107649, net125028,
         net112098, net112096, net112066, net112064, net110180, net99143,
         net99107, net99099, net83728, net83717, n96, net99193, net99127,
         net97350, net95120, net95119, net95115, net83707, net84368, net84360,
         net84337, net84335, net84310, net84309, net84299, net145688,
         net124986, net107667, n76, n77, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n90, n92, n94, n95, n98, n100, n101, n102, n103, n105,
         n106, n107, n116, n117, n119, n120, n121, n123, n124, n126, n127,
         n128, n130, n131, n132, n133, n134;
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U47 ( .A(n119), .B(n115), .ZN(SUM[22]) );
  NAND2_X1 U49 ( .A1(B[22]), .A2(A[22]), .ZN(n114) );
  NOR2_X1 U50 ( .A1(B[22]), .A2(A[22]), .ZN(n112) );
  XOR2_X1 U53 ( .A(net82621), .B(n118), .Z(SUM[21]) );
  XNOR2_X1 U56 ( .A(n123), .B(n122), .ZN(SUM[20]) );
  XOR2_X1 U62 ( .A(net112161), .B(n125), .Z(SUM[19]) );
  XNOR2_X1 U65 ( .A(net83718), .B(n129), .ZN(SUM[18]) );
  XNOR2_X1 U74 ( .A(net88223), .B(n136), .ZN(SUM[16]) );
  XNOR2_X1 U81 ( .A(n140), .B(n141), .ZN(SUM[15]) );
  AOI21_X1 U83 ( .B1(B[15]), .B2(net83123), .A(n116), .ZN(n140) );
  NOR2_X1 U75 ( .A1(net110243), .A2(net74518), .ZN(n136) );
  NAND2_X1 U82 ( .A1(net110231), .A2(A[14]), .ZN(n141) );
  XOR2_X1 U16 ( .A(net110231), .B(A[14]), .Z(SUM[14]) );
  NAND2_X1 U22 ( .A1(B[28]), .A2(A[28]), .ZN(n93) );
  NOR2_X1 U23 ( .A1(B[28]), .A2(A[28]), .ZN(n91) );
  XOR2_X1 U27 ( .A(B[27]), .B(A[27]), .Z(n97) );
  OAI21_X1 U19 ( .B1(net83728), .B2(n91), .A(n93), .ZN(n89) );
  NAND2_X1 U4 ( .A1(net107667), .A2(net83063), .ZN(net95089) );
  NAND2_X1 U5 ( .A1(net124986), .A2(net84368), .ZN(net84309) );
  NAND2_X1 U7 ( .A1(net84360), .A2(n76), .ZN(net84368) );
  OR2_X1 U8 ( .A1(net84337), .A2(net84329), .ZN(n76) );
  OR2_X1 U10 ( .A1(net84337), .A2(net145688), .ZN(net84360) );
  XOR2_X1 U15 ( .A(A[19]), .B(B[19]), .Z(n125) );
  NAND2_X1 U17 ( .A1(n117), .A2(n134), .ZN(net124986) );
  NAND2_X1 U18 ( .A1(n77), .A2(B[21]), .ZN(net84310) );
  INV_X1 U21 ( .A(A[21]), .ZN(net84335) );
  NAND2_X1 U24 ( .A1(A[19]), .A2(B[19]), .ZN(net84299) );
  NAND2_X1 U25 ( .A1(n117), .A2(n134), .ZN(net112161) );
  NAND2_X1 U26 ( .A1(net112066), .A2(net125028), .ZN(net124940) );
  XOR2_X1 U28 ( .A(A[21]), .B(B[21]), .Z(n118) );
  NAND2_X1 U29 ( .A1(B[21]), .A2(net84338), .ZN(net84337) );
  OAI21_X1 U30 ( .B1(net84303), .B2(net84299), .A(net84352), .ZN(net125026) );
  NAND2_X1 U32 ( .A1(net84349), .A2(n123), .ZN(net84350) );
  NAND2_X1 U33 ( .A1(net95119), .A2(n128), .ZN(net99193) );
  NAND2_X1 U34 ( .A1(net99193), .A2(A[27]), .ZN(net83717) );
  INV_X1 U37 ( .A(net97350), .ZN(n83) );
  OAI21_X1 U38 ( .B1(n133), .B2(net125031), .A(net95122), .ZN(net95119) );
  NAND2_X1 U39 ( .A1(net99127), .A2(n121), .ZN(net95120) );
  NAND2_X1 U40 ( .A1(net99158), .A2(net95120), .ZN(n82) );
  NAND2_X1 U52 ( .A1(n80), .A2(n81), .ZN(net116123) );
  NOR2_X1 U57 ( .A1(net99127), .A2(n124), .ZN(net99143) );
  NOR2_X1 U58 ( .A1(net99127), .A2(net99128), .ZN(net99126) );
  NAND2_X1 U59 ( .A1(net95115), .A2(net116113), .ZN(net97350) );
  NOR2_X1 U60 ( .A1(n82), .A2(net97350), .ZN(net99109) );
  NOR2_X1 U64 ( .A1(net83707), .A2(A[27]), .ZN(net116079) );
  NAND2_X1 U66 ( .A1(net116070), .A2(n79), .ZN(net95115) );
  XNOR2_X1 U71 ( .A(n131), .B(n126), .ZN(SUM[28]) );
  NAND2_X1 U76 ( .A1(n84), .A2(n85), .ZN(n96) );
  OR2_X1 U77 ( .A1(n124), .A2(net99107), .ZN(n85) );
  NAND2_X1 U79 ( .A1(net99099), .A2(net99143), .ZN(n84) );
  OAI21_X1 U84 ( .B1(net125031), .B2(net99050), .A(net95093), .ZN(net99099) );
  NAND2_X1 U89 ( .A1(net112096), .A2(net112093), .ZN(net112064) );
  INV_X1 U90 ( .A(net110228), .ZN(net112096) );
  INV_X1 U91 ( .A(net110245), .ZN(net110243) );
  NAND2_X1 U92 ( .A1(net110180), .A2(net112050), .ZN(net83718) );
  NAND2_X1 U93 ( .A1(net110228), .A2(net112050), .ZN(net84344) );
  INV_X1 U94 ( .A(n132), .ZN(net88213) );
  INV_X1 U97 ( .A(net110131), .ZN(net74518) );
  OAI21_X1 U98 ( .B1(net110243), .B2(net88223), .A(net110131), .ZN(net86108)
         );
  NAND2_X1 U100 ( .A1(net110228), .A2(net110223), .ZN(net110180) );
  AOI22_X1 U102 ( .A1(net124940), .A2(net125015), .B1(net125026), .B2(A[21]), 
        .ZN(net107649) );
  INV_X1 U104 ( .A(net125007), .ZN(net125015) );
  AOI22_X1 U105 ( .A1(net124940), .A2(net125015), .B1(net125026), .B2(A[21]), 
        .ZN(net83063) );
  AOI22_X1 U106 ( .A1(net125015), .A2(net112161), .B1(net125026), .B2(A[21]), 
        .ZN(net124943) );
  NAND2_X1 U107 ( .A1(net124940), .A2(net84366), .ZN(net84298) );
  INV_X1 U108 ( .A(net116138), .ZN(net84303) );
  NAND2_X1 U110 ( .A1(A[15]), .A2(B[15]), .ZN(net110220) );
  NAND2_X1 U111 ( .A1(B[16]), .A2(A[16]), .ZN(net110131) );
  CLKBUF_X1 U112 ( .A(A[15]), .Z(net83123) );
  CLKBUF_X1 U114 ( .A(B[14]), .Z(net110231) );
  OR2_X1 U118 ( .A1(A[20]), .A2(B[20]), .ZN(net84338) );
  OR2_X1 U119 ( .A1(B[20]), .A2(A[20]), .ZN(net116138) );
  CLKBUF_X1 U120 ( .A(A[20]), .Z(n86) );
  NAND2_X1 U121 ( .A1(B[20]), .A2(n86), .ZN(net84349) );
  NAND2_X1 U122 ( .A1(B[20]), .A2(n86), .ZN(net84352) );
  OR2_X1 U127 ( .A1(net116155), .A2(net95224), .ZN(n87) );
  INV_X1 U128 ( .A(net95222), .ZN(net116155) );
  NAND2_X1 U129 ( .A1(net125041), .A2(net99137), .ZN(net116153) );
  OAI21_X1 U130 ( .B1(net125031), .B2(net99050), .A(net95122), .ZN(net99158)
         );
  NAND2_X1 U134 ( .A1(net95089), .A2(net95236), .ZN(n88) );
  NAND2_X1 U137 ( .A1(A[23]), .A2(B[23]), .ZN(net95098) );
  OR2_X1 U138 ( .A1(n92), .A2(n114), .ZN(net95234) );
  INV_X1 U139 ( .A(A[23]), .ZN(n92) );
  NAND2_X1 U142 ( .A1(net99183), .A2(n90), .ZN(net95128) );
  XOR2_X1 U144 ( .A(A[23]), .B(B[23]), .Z(n111) );
  NAND2_X1 U145 ( .A1(net112059), .A2(net112060), .ZN(net110245) );
  NAND2_X1 U146 ( .A1(n94), .A2(n95), .ZN(net112050) );
  INV_X1 U147 ( .A(A[17]), .ZN(n95) );
  NAND2_X1 U150 ( .A1(A[17]), .A2(B[17]), .ZN(net110228) );
  NAND2_X1 U151 ( .A1(A[18]), .A2(B[18]), .ZN(net112065) );
  XNOR2_X1 U153 ( .A(n89), .B(net82778), .ZN(SUM[29]) );
  XNOR2_X1 U154 ( .A(B[29]), .B(A[29]), .ZN(net82778) );
  XNOR2_X1 U156 ( .A(n107), .B(n98), .ZN(SUM[26]) );
  XNOR2_X1 U158 ( .A(net125034), .B(n120), .ZN(SUM[24]) );
  INV_X1 U160 ( .A(net97351), .ZN(net125034) );
  NAND2_X1 U161 ( .A1(net145688), .A2(net84329), .ZN(net84366) );
  NAND2_X1 U162 ( .A1(net83063), .A2(net99137), .ZN(net99183) );
  NAND2_X1 U164 ( .A1(net112169), .A2(net99137), .ZN(net112166) );
  INV_X1 U166 ( .A(B[23]), .ZN(net95223) );
  OR2_X1 U167 ( .A1(net95223), .A2(n114), .ZN(net95222) );
  NOR2_X1 U170 ( .A1(n112), .A2(net95052), .ZN(n115) );
  NAND2_X1 U172 ( .A1(n100), .A2(n101), .ZN(net95093) );
  NAND2_X1 U174 ( .A1(A[25]), .A2(B[25]), .ZN(net116094) );
  XOR2_X1 U180 ( .A(A[25]), .B(B[25]), .Z(n104) );
  NAND2_X1 U182 ( .A1(A[24]), .A2(B[24]), .ZN(net116111) );
  NAND2_X1 U183 ( .A1(B[26]), .A2(A[26]), .ZN(net116113) );
  NAND2_X1 U184 ( .A1(n103), .A2(n102), .ZN(net116070) );
  OAI21_X1 U187 ( .B1(net116127), .B2(net116117), .A(n105), .ZN(n106) );
  NAND2_X1 U188 ( .A1(net116113), .A2(net116070), .ZN(n107) );
  NAND2_X1 U189 ( .A1(net112166), .A2(n87), .ZN(net112146) );
  INV_X1 U193 ( .A(n93), .ZN(net74529) );
  XNOR2_X1 U194 ( .A(net99109), .B(n97), .ZN(SUM[27]) );
  XNOR2_X1 U195 ( .A(n127), .B(n111), .ZN(SUM[23]) );
  INV_X1 U204 ( .A(B[27]), .ZN(net99106) );
  XNOR2_X1 U206 ( .A(net99126), .B(n104), .ZN(SUM[25]) );
  NOR2_X1 U212 ( .A1(net83123), .A2(B[15]), .ZN(n116) );
  NOR2_X1 U213 ( .A1(net88213), .A2(net84293), .ZN(n129) );
  NOR2_X1 U214 ( .A1(net84303), .A2(net84304), .ZN(n122) );
  XNOR2_X1 U216 ( .A(net86108), .B(net84344), .ZN(SUM[17]) );
  NAND4_X1 U2 ( .A1(net112098), .A2(net110245), .A3(net112050), .A4(n132), 
        .ZN(n117) );
  AND2_X1 U3 ( .A1(net124943), .A2(net99137), .ZN(n119) );
  NOR2_X1 U6 ( .A1(net116117), .A2(n130), .ZN(n120) );
  AND2_X1 U9 ( .A1(net116070), .A2(net116123), .ZN(n121) );
  AND2_X1 U11 ( .A1(net84298), .A2(net84299), .ZN(n123) );
  NOR2_X1 U12 ( .A1(net99106), .A2(net99092), .ZN(n124) );
  NOR2_X1 U13 ( .A1(n91), .A2(net74529), .ZN(n126) );
  AND2_X1 U14 ( .A1(net95128), .A2(n114), .ZN(n127) );
  AND2_X1 U20 ( .A1(net95120), .A2(n83), .ZN(n128) );
  AND2_X1 U31 ( .A1(B[24]), .A2(A[24]), .ZN(n130) );
  AND2_X1 U35 ( .A1(n96), .A2(net83717), .ZN(n131) );
  AND2_X1 U36 ( .A1(n96), .A2(net83717), .ZN(net83728) );
  OR2_X1 U41 ( .A1(B[18]), .A2(A[18]), .ZN(n132) );
  OR2_X1 U42 ( .A1(B[18]), .A2(A[18]), .ZN(net112093) );
  OAI211_X1 U43 ( .C1(net99166), .C2(net99082), .A(net95098), .B(net95234), 
        .ZN(n133) );
  OAI211_X1 U44 ( .C1(net99166), .C2(net99082), .A(net95098), .B(net95234), 
        .ZN(net99050) );
  NAND3_X1 U45 ( .A1(net97413), .A2(net112146), .A3(net95098), .ZN(net97351)
         );
  AND2_X1 U46 ( .A1(net112064), .A2(net112065), .ZN(n134) );
  AND2_X1 U48 ( .A1(net112064), .A2(net112065), .ZN(net125028) );
  OAI211_X1 U51 ( .C1(A[19]), .C2(B[19]), .A(A[21]), .B(net116138), .ZN(
        net125007) );
  OAI211_X1 U54 ( .C1(net84337), .C2(net84299), .A(net84349), .B(net84335), 
        .ZN(n77) );
  AND2_X1 U55 ( .A1(net116079), .A2(net95115), .ZN(net99092) );
  AND2_X1 U61 ( .A1(n88), .A2(net95234), .ZN(net97413) );
  AND2_X1 U63 ( .A1(net124943), .A2(net95222), .ZN(net112169) );
  INV_X1 U67 ( .A(net95093), .ZN(net116117) );
  OAI211_X1 U68 ( .C1(A[15]), .C2(B[15]), .A(B[14]), .B(A[14]), .ZN(net110221)
         );
  AND2_X1 U69 ( .A1(net84309), .A2(net84310), .ZN(net99137) );
  AND2_X1 U70 ( .A1(n90), .A2(B[23]), .ZN(net95224) );
  INV_X1 U72 ( .A(B[17]), .ZN(n94) );
  INV_X1 U73 ( .A(net86108), .ZN(net110223) );
  INV_X1 U78 ( .A(net116094), .ZN(n79) );
  INV_X1 U80 ( .A(n114), .ZN(net95052) );
  AND2_X1 U85 ( .A1(n106), .A2(net116123), .ZN(n98) );
  INV_X1 U86 ( .A(net116113), .ZN(net83707) );
  INV_X1 U87 ( .A(B[16]), .ZN(net112059) );
  INV_X1 U88 ( .A(A[16]), .ZN(net112060) );
  NAND4_X1 U95 ( .A1(net112098), .A2(net110245), .A3(net112050), .A4(n132), 
        .ZN(net112066) );
  NAND3_X1 U96 ( .A1(net110221), .A2(net110220), .A3(net110131), .ZN(net112098) );
  INV_X1 U99 ( .A(A[19]), .ZN(net145688) );
  INV_X1 U101 ( .A(B[19]), .ZN(net84329) );
  INV_X1 U103 ( .A(n112), .ZN(n90) );
  AND2_X1 U109 ( .A1(net84309), .A2(net84310), .ZN(net107667) );
  AND2_X1 U113 ( .A1(n90), .A2(A[23]), .ZN(net95236) );
  AND2_X1 U115 ( .A1(net110221), .A2(net110220), .ZN(net88223) );
  INV_X1 U116 ( .A(B[24]), .ZN(n101) );
  INV_X1 U117 ( .A(A[24]), .ZN(n100) );
  AND2_X1 U123 ( .A1(n121), .A2(B[27]), .ZN(net99107) );
  AND2_X1 U124 ( .A1(net95093), .A2(n121), .ZN(net95122) );
  INV_X1 U125 ( .A(net95236), .ZN(net99082) );
  AND2_X1 U126 ( .A1(net107667), .A2(net107649), .ZN(net99166) );
  AND2_X1 U131 ( .A1(net116153), .A2(n87), .ZN(net125031) );
  AND2_X1 U132 ( .A1(net107649), .A2(net95222), .ZN(net125041) );
  INV_X1 U133 ( .A(net112065), .ZN(net84293) );
  INV_X1 U135 ( .A(net84352), .ZN(net84304) );
  AND2_X1 U136 ( .A1(net116138), .A2(net84350), .ZN(net82621) );
  AND2_X1 U140 ( .A1(net97351), .A2(net95093), .ZN(net99128) );
  INV_X1 U141 ( .A(net116111), .ZN(net99127) );
  INV_X1 U143 ( .A(B[26]), .ZN(n103) );
  INV_X1 U148 ( .A(A[26]), .ZN(n102) );
  INV_X1 U149 ( .A(B[25]), .ZN(n80) );
  INV_X1 U152 ( .A(A[25]), .ZN(n81) );
  AND3_X1 U155 ( .A1(net112146), .A2(net95098), .A3(net97413), .ZN(net116127)
         );
  AND2_X1 U157 ( .A1(net116094), .A2(net116111), .ZN(n105) );
endmodule


module ALU_N32_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] , \ab[12][13] ,
         \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] , \ab[11][14] ,
         \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][12] ,
         \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] ,
         \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] ,
         \ab[8][0] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][15] , \ab[5][14] ,
         \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] ,
         \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][15] ,
         \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] ,
         \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] ,
         \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][8] , \ab[3][7] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][9] , \ab[2][8] ,
         \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] ,
         \ab[2][0] , \ab[1][15] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][1] , \ab[1][0] , \ab[0][15] , \ab[0][14] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][0] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[15][15] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][1] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][1] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , QA, QB,
         \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] ,
         \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] ,
         \A2[14] , n3, n4, n5, n6, n9, n11, n12, n15, n16, n17, n18, n19, n20,
         n21, n25, n26, n28, n29, n30, n31, n34, n36, n37, n38, n39, n40, n41,
         n49, n50, n51, n52, n53, n54, n62, n63, n99, n61, n60, n59, n58, n57,
         n56, n55, n48, n47, n46, n45, n44, n43, n42, n32, net74486, net74499,
         net76821, net76827, net76831, net76866, net76865, net76873, net76872,
         net77238, net82646, net82644, net82656, net82664, net82665, net82786,
         net82807, net82848, net82868, net82866, net83036, net83034, net83044,
         net83042, net83056, net83054, net83077, net83091, net83154, net83153,
         net83231, net83230, net83284, net83313, net83346, net83407, net83415,
         net83413, net83494, net83506, net83624, net83786, net86087, net86102,
         net86104, net88197, net88201, net88235, net88254, net94668, net95229,
         net99186, net110260, net112156, net95160, net83610, net74496,
         \ab[0][12] , net97393, net94632, \ab[3][9] , \ab[2][10] , net83140,
         net110254, ZA, net74508, net86070, \ab[4][9] , \SUMB[3][10] ,
         \SUMB[11][2] , \CARRYB[9][4] , \CARRYB[8][5] , \CARRYB[7][6] ,
         \CARRYB[6][7] , \CARRYB[5][8] , \CARRYB[4][9] , \CARRYB[11][2] ,
         \CARRYB[10][3] , net95231, n7, n23, \SUMB[9][4] , \SUMB[8][5] ,
         \SUMB[7][6] , \SUMB[6][7] , \SUMB[5][8] , \SUMB[4][9] , \SUMB[2][10] ,
         \SUMB[10][3] , \SUMB[10][2] , \CARRYB[9][3] , \CARRYB[8][4] ,
         \CARRYB[7][5] , \CARRYB[6][6] , \CARRYB[5][7] , \CARRYB[4][8] ,
         \CARRYB[3][9] , \CARRYB[2][10] , \CARRYB[10][2] , net97340, net83498,
         net83048, net82901, n10, \SUMB[9][3] , \SUMB[9][2] , \SUMB[8][4] ,
         \SUMB[7][5] , \SUMB[6][6] , \SUMB[5][7] , \SUMB[4][8] , \SUMB[3][9] ,
         \SUMB[2][9] , \CARRYB[9][2] , \CARRYB[8][3] , \CARRYB[7][4] ,
         \CARRYB[6][5] , \CARRYB[5][6] , \CARRYB[4][7] , \CARRYB[3][8] ,
         \CARRYB[2][9] , net83534, net82934, n8, n24, \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[7][4] , \SUMB[6][5] , \SUMB[5][6] , \SUMB[4][7] ,
         \SUMB[3][8] , \SUMB[2][8] , \CARRYB[8][2] , \CARRYB[7][3] ,
         \CARRYB[6][4] , \CARRYB[5][5] , \CARRYB[4][6] , \CARRYB[3][7] ,
         \CARRYB[2][8] , \SUMB[7][3] , \SUMB[7][2] , \CARRYB[7][2] , net83058,
         net82676, \ab[1][8] , \ab[0][9] , \ab[0][8] , \SUMB[6][4] ,
         \SUMB[6][3] , \CARRYB[6][3] , \SUMB[5][5] , \SUMB[5][4] ,
         \CARRYB[5][4] , \SUMB[4][6] , \SUMB[4][5] , \CARRYB[4][5] , net82974,
         \ab[8][6] , \SUMB[8][6] , \SUMB[7][7] , \CARRYB[9][5] ,
         \CARRYB[8][6] , net74503, n27, n22, n14, n13, \ab[3][6] , \ab[2][7] ,
         \ab[2][6] , \ab[1][7] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[2][7] ,
         \SUMB[2][6] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[2][7] ,
         \CARRYB[2][6] , net83003, net110253, net110252, \ab[13][2] ,
         \SUMB[9][5] , \SUMB[15][0] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][2] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[11][3] ,
         \SUMB[10][4] , \CARRYB[15][0] , \CARRYB[14][1] , \CARRYB[13][2] ,
         \CARRYB[13][1] , \CARRYB[12][2] , \CARRYB[11][3] , \CARRYB[10][4] ,
         n102, n103, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n125, n126, n127,
         n128, n129, n132, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n176, n177, n179, n180, n181, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n204, n205, n207, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n228, n229, n230, n231, n233, n234, n235, n236, n237, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n303, n306, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331;

  FA_X1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S14_15 ( .A(QA), .B(QB), .CI(\ab[15][15] ), .CO(\CARRYB[15][15] ), .S(
        \SUMB[15][15] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\CARRYB[13][8] ), .B(\ab[14][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_4 ( .A(\CARRYB[12][4] ), .B(\ab[13][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_8 ( .A(\CARRYB[12][8] ), .B(\ab[13][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\CARRYB[10][10] ), .B(\ab[11][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_7 ( .A(\CARRYB[8][7] ), .B(\ab[9][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\CARRYB[7][12] ), .B(\ab[8][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\CARRYB[6][1] ), .B(\ab[7][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_11 ( .A(\CARRYB[6][11] ), .B(\ab[7][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\CARRYB[6][12] ), .B(\ab[7][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\CARRYB[5][1] ), .B(\ab[6][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\CARRYB[5][2] ), .B(\ab[6][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_9 ( .A(\CARRYB[5][9] ), .B(\ab[6][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\SUMB[5][13] ), .B(\ab[6][12] ), .CI(\CARRYB[5][12] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\CARRYB[4][1] ), .B(\ab[5][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\CARRYB[4][2] ), .B(\ab[5][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_10 ( .A(\CARRYB[4][10] ), .B(\ab[5][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_12 ( .A(\CARRYB[4][12] ), .B(\ab[5][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\SUMB[4][14] ), .CI(\CARRYB[4][13] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\CARRYB[3][1] ), .B(\ab[4][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\CARRYB[3][2] ), .B(\ab[4][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\CARRYB[3][4] ), .B(\ab[4][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\CARRYB[3][11] ), .B(\ab[4][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\SUMB[3][14] ), .CI(\CARRYB[3][13] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_4 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n4), .CI(n20), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n6), .CI(n19), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n5), .CI(n18), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n3), .CI(n30), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(n16), .B(\ab[2][4] ), .CI(n29), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n11), .CI(n26), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S3_2_14 ( .A(n17), .B(\ab[2][14] ), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  XOR2_X1 U17 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(n18) );
  XOR2_X1 U18 ( .A(n323), .B(\ab[0][3] ), .Z(n19) );
  XOR2_X1 U19 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n20) );
  XOR2_X1 U27 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n28) );
  XOR2_X1 U28 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n29) );
  XOR2_X1 U32 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  XOR2_X1 U38 ( .A(\CARRYB[15][7] ), .B(\SUMB[15][8] ), .Z(n37) );
  XOR2_X1 U39 ( .A(\CARRYB[15][9] ), .B(\SUMB[15][10] ), .Z(n38) );
  XOR2_X1 U40 ( .A(\CARRYB[15][11] ), .B(\SUMB[15][12] ), .Z(n39) );
  XOR2_X1 U41 ( .A(\CARRYB[15][13] ), .B(\SUMB[15][14] ), .Z(n40) );
  XOR2_X1 U52 ( .A(\SUMB[15][7] ), .B(\CARRYB[15][6] ), .Z(n51) );
  XOR2_X1 U53 ( .A(\CARRYB[15][8] ), .B(\SUMB[15][9] ), .Z(n52) );
  XOR2_X1 U54 ( .A(\CARRYB[15][10] ), .B(\SUMB[15][11] ), .Z(n53) );
  XOR2_X1 U55 ( .A(\CARRYB[15][12] ), .B(\SUMB[15][13] ), .Z(n54) );
  XOR2_X1 U63 ( .A(\CARRYB[15][14] ), .B(\SUMB[15][15] ), .Z(n62) );
  NOR2_X1 U98 ( .A1(n314), .A2(net83036), .ZN(\ab[9][9] ) );
  NOR2_X1 U99 ( .A1(n314), .A2(net83624), .ZN(\ab[9][8] ) );
  NOR2_X1 U100 ( .A1(n314), .A2(net83313), .ZN(\ab[9][7] ) );
  NOR2_X1 U101 ( .A1(n314), .A2(net83346), .ZN(\ab[9][6] ) );
  NOR2_X1 U102 ( .A1(n314), .A2(n318), .ZN(\ab[9][5] ) );
  NOR2_X1 U103 ( .A1(n314), .A2(n303), .ZN(\ab[9][4] ) );
  NOR2_X1 U104 ( .A1(n314), .A2(n306), .ZN(\ab[9][3] ) );
  NOR2_X1 U105 ( .A1(n314), .A2(net74486), .ZN(\ab[9][2] ) );
  NOR2_X1 U106 ( .A1(n314), .A2(n132), .ZN(\ab[9][1] ) );
  NOR2_X1 U108 ( .A1(n314), .A2(net83506), .ZN(\ab[9][14] ) );
  NOR2_X1 U109 ( .A1(n314), .A2(net83154), .ZN(\ab[9][13] ) );
  NOR2_X1 U110 ( .A1(n314), .A2(net83415), .ZN(\ab[9][12] ) );
  NOR2_X1 U111 ( .A1(n314), .A2(net82848), .ZN(\ab[9][11] ) );
  NOR2_X1 U112 ( .A1(n314), .A2(net95229), .ZN(\ab[9][10] ) );
  NOR2_X1 U113 ( .A1(n314), .A2(n322), .ZN(\ab[9][0] ) );
  NOR2_X1 U114 ( .A1(net83036), .A2(net74508), .ZN(\ab[8][9] ) );
  NOR2_X1 U115 ( .A1(net83624), .A2(net74508), .ZN(\ab[8][8] ) );
  NOR2_X1 U116 ( .A1(net83313), .A2(net74508), .ZN(\ab[8][7] ) );
  NOR2_X1 U118 ( .A1(n201), .A2(net74508), .ZN(\ab[8][5] ) );
  NOR2_X1 U119 ( .A1(n303), .A2(net74508), .ZN(\ab[8][4] ) );
  NOR2_X1 U120 ( .A1(n306), .A2(net74508), .ZN(\ab[8][3] ) );
  NOR2_X1 U121 ( .A1(net74486), .A2(net74508), .ZN(\ab[8][2] ) );
  NOR2_X1 U122 ( .A1(n132), .A2(net74508), .ZN(\ab[8][1] ) );
  NOR2_X1 U124 ( .A1(net83506), .A2(net74508), .ZN(\ab[8][14] ) );
  NOR2_X1 U125 ( .A1(net83154), .A2(net74508), .ZN(\ab[8][13] ) );
  NOR2_X1 U126 ( .A1(net83415), .A2(net74508), .ZN(\ab[8][12] ) );
  NOR2_X1 U127 ( .A1(net82848), .A2(net74508), .ZN(\ab[8][11] ) );
  NOR2_X1 U128 ( .A1(net95229), .A2(net74508), .ZN(\ab[8][10] ) );
  NOR2_X1 U129 ( .A1(n322), .A2(net74508), .ZN(\ab[8][0] ) );
  NOR2_X1 U130 ( .A1(net83036), .A2(n315), .ZN(\ab[7][9] ) );
  NOR2_X1 U131 ( .A1(net83624), .A2(n315), .ZN(\ab[7][8] ) );
  NOR2_X1 U132 ( .A1(net83313), .A2(n315), .ZN(\ab[7][7] ) );
  NOR2_X1 U133 ( .A1(net83346), .A2(n315), .ZN(\ab[7][6] ) );
  NOR2_X1 U134 ( .A1(n201), .A2(n315), .ZN(\ab[7][5] ) );
  NOR2_X1 U135 ( .A1(n303), .A2(n315), .ZN(\ab[7][4] ) );
  NOR2_X1 U136 ( .A1(n306), .A2(n315), .ZN(\ab[7][3] ) );
  NOR2_X1 U137 ( .A1(net74486), .A2(n315), .ZN(\ab[7][2] ) );
  NOR2_X1 U138 ( .A1(n132), .A2(n315), .ZN(\ab[7][1] ) );
  NOR2_X1 U140 ( .A1(net83506), .A2(n315), .ZN(\ab[7][14] ) );
  NOR2_X1 U141 ( .A1(net83154), .A2(n315), .ZN(\ab[7][13] ) );
  NOR2_X1 U142 ( .A1(net83415), .A2(n315), .ZN(\ab[7][12] ) );
  NOR2_X1 U143 ( .A1(net82848), .A2(n315), .ZN(\ab[7][11] ) );
  NOR2_X1 U144 ( .A1(net83048), .A2(n315), .ZN(\ab[7][10] ) );
  NOR2_X1 U145 ( .A1(n322), .A2(n315), .ZN(\ab[7][0] ) );
  NOR2_X1 U146 ( .A1(net83036), .A2(n316), .ZN(\ab[6][9] ) );
  NOR2_X1 U147 ( .A1(net83624), .A2(n316), .ZN(\ab[6][8] ) );
  NOR2_X1 U148 ( .A1(net83313), .A2(n316), .ZN(\ab[6][7] ) );
  NOR2_X1 U149 ( .A1(net83346), .A2(n316), .ZN(\ab[6][6] ) );
  NOR2_X1 U150 ( .A1(n201), .A2(n316), .ZN(\ab[6][5] ) );
  NOR2_X1 U151 ( .A1(n303), .A2(n316), .ZN(\ab[6][4] ) );
  NOR2_X1 U152 ( .A1(n306), .A2(n316), .ZN(\ab[6][3] ) );
  NOR2_X1 U153 ( .A1(net74486), .A2(n316), .ZN(\ab[6][2] ) );
  NOR2_X1 U154 ( .A1(n132), .A2(n316), .ZN(\ab[6][1] ) );
  NOR2_X1 U156 ( .A1(net83506), .A2(n316), .ZN(\ab[6][14] ) );
  NOR2_X1 U157 ( .A1(net83154), .A2(n316), .ZN(\ab[6][13] ) );
  NOR2_X1 U158 ( .A1(net83415), .A2(n316), .ZN(\ab[6][12] ) );
  NOR2_X1 U159 ( .A1(net82848), .A2(n316), .ZN(\ab[6][11] ) );
  NOR2_X1 U160 ( .A1(net83048), .A2(n316), .ZN(\ab[6][10] ) );
  NOR2_X1 U161 ( .A1(n322), .A2(n316), .ZN(\ab[6][0] ) );
  NOR2_X1 U162 ( .A1(net83036), .A2(n317), .ZN(\ab[5][9] ) );
  NOR2_X1 U163 ( .A1(net83624), .A2(n317), .ZN(\ab[5][8] ) );
  NOR2_X1 U164 ( .A1(net83313), .A2(n317), .ZN(\ab[5][7] ) );
  NOR2_X1 U165 ( .A1(net83346), .A2(n317), .ZN(\ab[5][6] ) );
  NOR2_X1 U166 ( .A1(n318), .A2(n317), .ZN(\ab[5][5] ) );
  NOR2_X1 U167 ( .A1(n303), .A2(n317), .ZN(\ab[5][4] ) );
  NOR2_X1 U168 ( .A1(n306), .A2(n317), .ZN(\ab[5][3] ) );
  NOR2_X1 U169 ( .A1(net74486), .A2(n317), .ZN(\ab[5][2] ) );
  NOR2_X1 U170 ( .A1(n132), .A2(n317), .ZN(\ab[5][1] ) );
  NOR2_X1 U172 ( .A1(net83506), .A2(n317), .ZN(\ab[5][14] ) );
  NOR2_X1 U173 ( .A1(net83154), .A2(n317), .ZN(\ab[5][13] ) );
  NOR2_X1 U174 ( .A1(net83415), .A2(n317), .ZN(\ab[5][12] ) );
  NOR2_X1 U175 ( .A1(net82848), .A2(n317), .ZN(\ab[5][11] ) );
  NOR2_X1 U176 ( .A1(net83048), .A2(n317), .ZN(\ab[5][10] ) );
  NOR2_X1 U177 ( .A1(n322), .A2(n317), .ZN(\ab[5][0] ) );
  NOR2_X1 U179 ( .A1(net83624), .A2(net76873), .ZN(\ab[4][8] ) );
  NOR2_X1 U180 ( .A1(net83313), .A2(net76872), .ZN(\ab[4][7] ) );
  NOR2_X1 U181 ( .A1(net83346), .A2(net76873), .ZN(\ab[4][6] ) );
  NOR2_X1 U182 ( .A1(n201), .A2(net76872), .ZN(\ab[4][5] ) );
  NOR2_X1 U183 ( .A1(n303), .A2(net76873), .ZN(\ab[4][4] ) );
  NOR2_X1 U184 ( .A1(n306), .A2(net76872), .ZN(\ab[4][3] ) );
  NOR2_X1 U185 ( .A1(net74486), .A2(net76873), .ZN(\ab[4][2] ) );
  NOR2_X1 U186 ( .A1(n132), .A2(net76872), .ZN(\ab[4][1] ) );
  NOR2_X1 U188 ( .A1(net83506), .A2(net76873), .ZN(\ab[4][14] ) );
  NOR2_X1 U189 ( .A1(net83154), .A2(net76872), .ZN(\ab[4][13] ) );
  NOR2_X1 U190 ( .A1(net83415), .A2(net76873), .ZN(\ab[4][12] ) );
  NOR2_X1 U191 ( .A1(net82848), .A2(net76872), .ZN(\ab[4][11] ) );
  NOR2_X1 U192 ( .A1(net83048), .A2(net76872), .ZN(\ab[4][10] ) );
  NOR2_X1 U193 ( .A1(n322), .A2(net76872), .ZN(\ab[4][0] ) );
  NOR2_X1 U195 ( .A1(net83624), .A2(net76866), .ZN(\ab[3][8] ) );
  NOR2_X1 U196 ( .A1(net83313), .A2(net76866), .ZN(\ab[3][7] ) );
  NOR2_X1 U198 ( .A1(n201), .A2(net76866), .ZN(\ab[3][5] ) );
  NOR2_X1 U199 ( .A1(n303), .A2(net74503), .ZN(\ab[3][4] ) );
  NOR2_X1 U200 ( .A1(n306), .A2(net76866), .ZN(\ab[3][3] ) );
  NOR2_X1 U201 ( .A1(net74486), .A2(net74503), .ZN(\ab[3][2] ) );
  NOR2_X1 U202 ( .A1(n132), .A2(net76866), .ZN(\ab[3][1] ) );
  NOR2_X1 U204 ( .A1(net83506), .A2(net76866), .ZN(\ab[3][14] ) );
  NOR2_X1 U205 ( .A1(net86104), .A2(net76866), .ZN(\ab[3][13] ) );
  NOR2_X1 U206 ( .A1(net83415), .A2(net76865), .ZN(\ab[3][12] ) );
  NOR2_X1 U207 ( .A1(net82848), .A2(net76865), .ZN(\ab[3][11] ) );
  NOR2_X1 U208 ( .A1(net83048), .A2(net76865), .ZN(\ab[3][10] ) );
  NOR2_X1 U209 ( .A1(n322), .A2(net76866), .ZN(\ab[3][0] ) );
  NOR2_X1 U211 ( .A1(net99186), .A2(net97393), .ZN(\ab[2][8] ) );
  NOR2_X1 U214 ( .A1(n201), .A2(net97393), .ZN(\ab[2][5] ) );
  NOR2_X1 U215 ( .A1(n319), .A2(net83786), .ZN(\ab[2][4] ) );
  NOR2_X1 U216 ( .A1(n320), .A2(net83786), .ZN(\ab[2][3] ) );
  NOR2_X1 U217 ( .A1(net74486), .A2(net83786), .ZN(\ab[2][2] ) );
  NOR2_X1 U218 ( .A1(n132), .A2(net83786), .ZN(\ab[2][1] ) );
  NOR2_X1 U220 ( .A1(net83506), .A2(net97393), .ZN(\ab[2][14] ) );
  NOR2_X1 U221 ( .A1(net86104), .A2(net97393), .ZN(\ab[2][13] ) );
  NOR2_X1 U222 ( .A1(net82807), .A2(net97393), .ZN(\ab[2][12] ) );
  NOR2_X1 U225 ( .A1(n322), .A2(net83786), .ZN(\ab[2][0] ) );
  NOR2_X1 U230 ( .A1(n318), .A2(net83230), .ZN(\ab[1][5] ) );
  NOR2_X1 U231 ( .A1(n319), .A2(net83230), .ZN(\ab[1][4] ) );
  NOR2_X1 U232 ( .A1(n320), .A2(net83230), .ZN(\ab[1][3] ) );
  NOR2_X1 U234 ( .A1(n132), .A2(net83231), .ZN(\ab[1][1] ) );
  NOR2_X1 U241 ( .A1(n322), .A2(net83230), .ZN(\ab[1][0] ) );
  NOR2_X1 U259 ( .A1(net83036), .A2(n310), .ZN(\ab[14][9] ) );
  NOR2_X1 U260 ( .A1(net83624), .A2(n310), .ZN(\ab[14][8] ) );
  NOR2_X1 U261 ( .A1(net83313), .A2(n310), .ZN(\ab[14][7] ) );
  NOR2_X1 U262 ( .A1(net83346), .A2(n310), .ZN(\ab[14][6] ) );
  NOR2_X1 U263 ( .A1(n318), .A2(n310), .ZN(\ab[14][5] ) );
  NOR2_X1 U264 ( .A1(n303), .A2(n310), .ZN(\ab[14][4] ) );
  NOR2_X1 U265 ( .A1(n306), .A2(n310), .ZN(\ab[14][3] ) );
  NOR2_X1 U266 ( .A1(net74486), .A2(n310), .ZN(\ab[14][2] ) );
  NOR2_X1 U267 ( .A1(n132), .A2(n310), .ZN(\ab[14][1] ) );
  NOR2_X1 U269 ( .A1(net83506), .A2(n310), .ZN(\ab[14][14] ) );
  NOR2_X1 U270 ( .A1(net83154), .A2(n310), .ZN(\ab[14][13] ) );
  NOR2_X1 U271 ( .A1(net83415), .A2(n310), .ZN(\ab[14][12] ) );
  NOR2_X1 U272 ( .A1(net82848), .A2(n310), .ZN(\ab[14][11] ) );
  NOR2_X1 U273 ( .A1(net95229), .A2(n310), .ZN(\ab[14][10] ) );
  NOR2_X1 U274 ( .A1(n322), .A2(n310), .ZN(\ab[14][0] ) );
  NOR2_X1 U275 ( .A1(net83036), .A2(n102), .ZN(\ab[13][9] ) );
  NOR2_X1 U276 ( .A1(net83624), .A2(n102), .ZN(\ab[13][8] ) );
  NOR2_X1 U277 ( .A1(net83313), .A2(n102), .ZN(\ab[13][7] ) );
  NOR2_X1 U278 ( .A1(net83346), .A2(n102), .ZN(\ab[13][6] ) );
  NOR2_X1 U279 ( .A1(n201), .A2(n102), .ZN(\ab[13][5] ) );
  NOR2_X1 U280 ( .A1(n303), .A2(n102), .ZN(\ab[13][4] ) );
  NOR2_X1 U281 ( .A1(n306), .A2(n102), .ZN(\ab[13][3] ) );
  NOR2_X1 U283 ( .A1(n132), .A2(n102), .ZN(\ab[13][1] ) );
  NOR2_X1 U285 ( .A1(net83506), .A2(n102), .ZN(\ab[13][14] ) );
  NOR2_X1 U286 ( .A1(net83154), .A2(n102), .ZN(\ab[13][13] ) );
  NOR2_X1 U287 ( .A1(net83415), .A2(n102), .ZN(\ab[13][12] ) );
  NOR2_X1 U288 ( .A1(net82848), .A2(n102), .ZN(\ab[13][11] ) );
  NOR2_X1 U289 ( .A1(net95229), .A2(n102), .ZN(\ab[13][10] ) );
  NOR2_X1 U290 ( .A1(n322), .A2(n102), .ZN(\ab[13][0] ) );
  NOR2_X1 U291 ( .A1(net83036), .A2(n311), .ZN(\ab[12][9] ) );
  NOR2_X1 U292 ( .A1(net83624), .A2(n311), .ZN(\ab[12][8] ) );
  NOR2_X1 U293 ( .A1(net83313), .A2(n311), .ZN(\ab[12][7] ) );
  NOR2_X1 U294 ( .A1(net83346), .A2(n311), .ZN(\ab[12][6] ) );
  NOR2_X1 U295 ( .A1(n201), .A2(n311), .ZN(\ab[12][5] ) );
  NOR2_X1 U296 ( .A1(n303), .A2(n311), .ZN(\ab[12][4] ) );
  NOR2_X1 U297 ( .A1(n320), .A2(n311), .ZN(\ab[12][3] ) );
  NOR2_X1 U298 ( .A1(net74486), .A2(n311), .ZN(\ab[12][2] ) );
  NOR2_X1 U299 ( .A1(n132), .A2(n311), .ZN(\ab[12][1] ) );
  NOR2_X1 U301 ( .A1(net83506), .A2(n311), .ZN(\ab[12][14] ) );
  NOR2_X1 U302 ( .A1(net83154), .A2(n311), .ZN(\ab[12][13] ) );
  NOR2_X1 U303 ( .A1(net83415), .A2(n311), .ZN(\ab[12][12] ) );
  NOR2_X1 U304 ( .A1(net82848), .A2(n311), .ZN(\ab[12][11] ) );
  NOR2_X1 U305 ( .A1(net95229), .A2(n311), .ZN(\ab[12][10] ) );
  NOR2_X1 U306 ( .A1(n322), .A2(n311), .ZN(\ab[12][0] ) );
  NOR2_X1 U307 ( .A1(net83036), .A2(n312), .ZN(\ab[11][9] ) );
  NOR2_X1 U308 ( .A1(net83624), .A2(n312), .ZN(\ab[11][8] ) );
  NOR2_X1 U309 ( .A1(net83313), .A2(n312), .ZN(\ab[11][7] ) );
  NOR2_X1 U310 ( .A1(net83346), .A2(n312), .ZN(\ab[11][6] ) );
  NOR2_X1 U311 ( .A1(n201), .A2(n312), .ZN(\ab[11][5] ) );
  NOR2_X1 U312 ( .A1(n303), .A2(n312), .ZN(\ab[11][4] ) );
  NOR2_X1 U313 ( .A1(n306), .A2(n312), .ZN(\ab[11][3] ) );
  NOR2_X1 U314 ( .A1(net74486), .A2(n312), .ZN(\ab[11][2] ) );
  NOR2_X1 U315 ( .A1(n132), .A2(n312), .ZN(\ab[11][1] ) );
  NOR2_X1 U317 ( .A1(net83506), .A2(n312), .ZN(\ab[11][14] ) );
  NOR2_X1 U318 ( .A1(net83154), .A2(n312), .ZN(\ab[11][13] ) );
  NOR2_X1 U319 ( .A1(net83415), .A2(n312), .ZN(\ab[11][12] ) );
  NOR2_X1 U320 ( .A1(net82848), .A2(n312), .ZN(\ab[11][11] ) );
  NOR2_X1 U321 ( .A1(net95229), .A2(n312), .ZN(\ab[11][10] ) );
  NOR2_X1 U322 ( .A1(n322), .A2(n312), .ZN(\ab[11][0] ) );
  NOR2_X1 U323 ( .A1(net83036), .A2(n313), .ZN(\ab[10][9] ) );
  NOR2_X1 U324 ( .A1(net83624), .A2(n313), .ZN(\ab[10][8] ) );
  NOR2_X1 U325 ( .A1(net83313), .A2(n313), .ZN(\ab[10][7] ) );
  NOR2_X1 U326 ( .A1(net83346), .A2(n313), .ZN(\ab[10][6] ) );
  NOR2_X1 U327 ( .A1(n201), .A2(n313), .ZN(\ab[10][5] ) );
  NOR2_X1 U328 ( .A1(n303), .A2(n313), .ZN(\ab[10][4] ) );
  NOR2_X1 U329 ( .A1(n306), .A2(n313), .ZN(\ab[10][3] ) );
  NOR2_X1 U330 ( .A1(net74486), .A2(n313), .ZN(\ab[10][2] ) );
  NOR2_X1 U331 ( .A1(n132), .A2(n313), .ZN(\ab[10][1] ) );
  NOR2_X1 U333 ( .A1(net83506), .A2(n313), .ZN(\ab[10][14] ) );
  NOR2_X1 U334 ( .A1(net83154), .A2(n313), .ZN(\ab[10][13] ) );
  NOR2_X1 U335 ( .A1(net83415), .A2(n313), .ZN(\ab[10][12] ) );
  NOR2_X1 U336 ( .A1(net82848), .A2(n313), .ZN(\ab[10][11] ) );
  NOR2_X1 U337 ( .A1(net95229), .A2(n313), .ZN(\ab[10][10] ) );
  NOR2_X1 U338 ( .A1(n322), .A2(n313), .ZN(\ab[10][0] ) );
  NOR2_X1 U343 ( .A1(n318), .A2(net83494), .ZN(\ab[0][5] ) );
  NOR2_X1 U344 ( .A1(n319), .A2(net83494), .ZN(\ab[0][4] ) );
  NOR2_X1 U345 ( .A1(n320), .A2(net83494), .ZN(\ab[0][3] ) );
  NOR2_X1 U346 ( .A1(net74486), .A2(net82901), .ZN(\ab[0][2] ) );
  NOR2_X1 U347 ( .A1(n132), .A2(net83494), .ZN(\ab[0][1] ) );
  NOR2_X1 U357 ( .A1(n322), .A2(net88254), .ZN(PRODUCT[0]) );
  NOR2_X1 U194 ( .A1(net83036), .A2(net76866), .ZN(\ab[3][9] ) );
  NOR2_X1 U223 ( .A1(net94632), .A2(net97393), .ZN(\ab[2][11] ) );
  NOR2_X1 U251 ( .A1(net83407), .A2(n110), .ZN(\ab[15][15] ) );
  XOR2_X1 U97 ( .A(\CARRYB[15][15] ), .B(n111), .Z(n63) );
  NOR2_X1 U258 ( .A1(n110), .A2(n111), .ZN(n99) );
  NOR2_X1 U355 ( .A1(net82665), .A2(n109), .ZN(QB) );
  NOR2_X1 U356 ( .A1(A[15]), .A2(n109), .ZN(QA) );
  NOR2_X1 U34 ( .A1(n110), .A2(n109), .ZN(ZA) );
  NOR2_X1 U178 ( .A1(net83036), .A2(net76872), .ZN(\ab[4][9] ) );
  FA_X1 S2_12_1 ( .A(\CARRYB[11][1] ), .B(\ab[12][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n7), .CI(n23), .CO(\CARRYB[2][10] ), .S(
        \SUMB[2][10] ) );
  FA_X1 S2_4_9 ( .A(\CARRYB[3][9] ), .B(\ab[4][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_5_8 ( .A(\CARRYB[4][8] ), .B(\ab[5][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_6_7 ( .A(\CARRYB[5][7] ), .B(\ab[6][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_7_6 ( .A(\CARRYB[6][6] ), .B(\ab[7][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_8_5 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_9_4 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_10_3 ( .A(\CARRYB[9][3] ), .B(\ab[10][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_11_1 ( .A(\CARRYB[10][1] ), .B(\ab[11][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\CARRYB[10][2] ), .B(\ab[11][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  NOR2_X1 U352 ( .A1(net74496), .A2(net82901), .ZN(\ab[0][12] ) );
  NOR2_X1 U224 ( .A1(net97393), .A2(net83048), .ZN(\ab[2][10] ) );
  FA_X1 S2_3_9 ( .A(\CARRYB[2][9] ), .B(\ab[3][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n21), .CI(n10), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_4_8 ( .A(\CARRYB[3][8] ), .B(\ab[4][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_5_7 ( .A(\CARRYB[4][7] ), .B(\ab[5][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_6_6 ( .A(\CARRYB[5][6] ), .B(\ab[6][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_7_5 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_8_4 ( .A(\CARRYB[7][4] ), .B(\ab[8][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_9_3 ( .A(\CARRYB[8][3] ), .B(\ab[9][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_10_1 ( .A(\CARRYB[9][1] ), .B(\ab[10][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\CARRYB[9][2] ), .B(\ab[10][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n8), .CI(n24), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_4_7 ( .A(\CARRYB[3][7] ), .B(\ab[4][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_5_6 ( .A(\CARRYB[4][6] ), .B(\ab[5][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_6_5 ( .A(\CARRYB[5][5] ), .B(\ab[6][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_7_4 ( .A(\CARRYB[6][4] ), .B(\ab[7][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_8_3 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_9_1 ( .A(\CARRYB[8][1] ), .B(\ab[9][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\CARRYB[8][2] ), .B(\ab[9][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_8_1 ( .A(\CARRYB[7][1] ), .B(\ab[8][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\CARRYB[7][2] ), .B(\ab[8][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  NOR2_X1 U339 ( .A1(net82676), .A2(net88254), .ZN(\ab[0][9] ) );
  FA_X1 S2_7_2 ( .A(\CARRYB[6][2] ), .B(\ab[7][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\CARRYB[6][3] ), .B(\ab[7][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_6_3 ( .A(\CARRYB[5][3] ), .B(\ab[6][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\CARRYB[5][4] ), .B(\ab[6][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_5_4 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\CARRYB[4][5] ), .B(\ab[5][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  NOR2_X1 U117 ( .A1(net83346), .A2(net74508), .ZN(\ab[8][6] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_8_6 ( .A(\CARRYB[7][6] ), .B(\ab[8][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_3_5 ( .A(\CARRYB[2][5] ), .B(\ab[3][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n14), .CI(n27), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  NOR2_X1 U197 ( .A1(net83346), .A2(net76866), .ZN(\ab[3][6] ) );
  NOR2_X1 U212 ( .A1(n103), .A2(net83786), .ZN(\ab[2][7] ) );
  XOR2_X1 U21 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(n22) );
  FA_X1 S2_3_7 ( .A(\CARRYB[2][7] ), .B(\ab[3][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n13), .CI(n22), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_4_5 ( .A(\CARRYB[3][5] ), .B(\ab[4][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\CARRYB[3][6] ), .B(\ab[4][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_3_6 ( .A(\CARRYB[2][6] ), .B(\ab[3][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_9_5 ( .A(\CARRYB[8][5] ), .B(\ab[9][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_10_4 ( .A(\CARRYB[9][4] ), .B(\ab[10][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_11_3 ( .A(\CARRYB[10][3] ), .B(\ab[11][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_13_1 ( .A(\CARRYB[12][1] ), .B(\ab[13][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_12_2 ( .A(\CARRYB[11][2] ), .B(\ab[12][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  NOR2_X1 U282 ( .A1(net74486), .A2(n102), .ZN(\ab[13][2] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_13_2 ( .A(\CARRYB[12][2] ), .B(\ab[13][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_14_1 ( .A(\CARRYB[13][1] ), .B(\ab[14][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S4_0 ( .A(\CARRYB[14][0] ), .B(\ab[15][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  NAND2_X1 U6 ( .A1(\SUMB[15][0] ), .A2(net76831), .ZN(net110253) );
  NAND2_X1 U24 ( .A1(\SUMB[15][0] ), .A2(net76827), .ZN(net110252) );
  XNOR2_X1 U25 ( .A(net83003), .B(\SUMB[11][4] ), .ZN(\SUMB[12][3] ) );
  XNOR2_X1 U26 ( .A(\CARRYB[11][3] ), .B(\ab[12][3] ), .ZN(net83003) );
  INV_X1 U30 ( .A(A[13]), .ZN(n102) );
  INV_X2 U36 ( .A(B[2]), .ZN(net74486) );
  NAND2_X1 U37 ( .A1(\CARRYB[11][3] ), .A2(\ab[12][3] ), .ZN(net82646) );
  NAND2_X1 U42 ( .A1(\SUMB[11][4] ), .A2(\CARRYB[11][3] ), .ZN(net82644) );
  NAND2_X1 U50 ( .A1(\CARRYB[9][5] ), .A2(\ab[10][5] ), .ZN(net83044) );
  XNOR2_X1 U51 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .ZN(net83091) );
  INV_X1 U66 ( .A(net83284), .ZN(\ab[1][7] ) );
  INV_X1 U73 ( .A(B[7]), .ZN(net83313) );
  INV_X1 U74 ( .A(B[7]), .ZN(n103) );
  INV_X1 U76 ( .A(A[3]), .ZN(net74503) );
  CLKBUF_X3 U77 ( .A(net74503), .Z(net76866) );
  INV_X2 U79 ( .A(B[6]), .ZN(net83346) );
  XNOR2_X1 U83 ( .A(\ab[0][8] ), .B(net83284), .ZN(n27) );
  NAND2_X1 U84 ( .A1(\SUMB[9][6] ), .A2(\CARRYB[9][5] ), .ZN(net83042) );
  XNOR2_X1 U85 ( .A(net82974), .B(\SUMB[6][8] ), .ZN(\SUMB[7][7] ) );
  XNOR2_X1 U86 ( .A(\CARRYB[6][7] ), .B(\ab[7][7] ), .ZN(net82974) );
  CLKBUF_X1 U89 ( .A(net82901), .Z(net83494) );
  INV_X1 U90 ( .A(A[0]), .ZN(net83058) );
  INV_X1 U91 ( .A(net83058), .ZN(net82934) );
  INV_X1 U93 ( .A(B[9]), .ZN(net82676) );
  INV_X1 U94 ( .A(net82676), .ZN(net83034) );
  NOR2_X1 U210 ( .A1(net99186), .A2(net88254), .ZN(\ab[0][8] ) );
  NOR2_X1 U226 ( .A1(net86104), .A2(net88254), .ZN(net83153) );
  INV_X1 U227 ( .A(A[8]), .ZN(net74508) );
  XNOR2_X1 U229 ( .A(net97340), .B(net83534), .ZN(n24) );
  NAND2_X1 U233 ( .A1(B[10]), .A2(net82934), .ZN(net83534) );
  NAND2_X1 U236 ( .A1(net82934), .A2(net95160), .ZN(net95231) );
  INV_X1 U340 ( .A(A[1]), .ZN(net83231) );
  NOR2_X1 U342 ( .A1(net82676), .A2(net83231), .ZN(net97340) );
  NOR2_X1 U349 ( .A1(net82901), .A2(net83048), .ZN(net83498) );
  INV_X1 U350 ( .A(B[10]), .ZN(net83048) );
  INV_X1 U354 ( .A(A[0]), .ZN(net82901) );
  NOR2_X1 U358 ( .A1(net94632), .A2(net82901), .ZN(net83610) );
  XNOR2_X1 U360 ( .A(\CARRYB[2][10] ), .B(\ab[3][10] ), .ZN(net86070) );
  XNOR2_X1 U361 ( .A(\ab[0][12] ), .B(n107), .ZN(n23) );
  NAND2_X1 U362 ( .A1(B[11]), .A2(A[1]), .ZN(n107) );
  NOR2_X1 U363 ( .A1(net94632), .A2(net95231), .ZN(n7) );
  NAND2_X1 U365 ( .A1(\CARRYB[6][7] ), .A2(\ab[7][7] ), .ZN(net82664) );
  XNOR2_X1 U366 ( .A(\CARRYB[5][8] ), .B(\ab[6][8] ), .ZN(net83077) );
  NAND2_X1 U367 ( .A1(\CARRYB[5][8] ), .A2(\ab[6][8] ), .ZN(net82868) );
  NAND2_X1 U368 ( .A1(\SUMB[5][9] ), .A2(\CARRYB[5][8] ), .ZN(net82866) );
  XNOR2_X1 U369 ( .A(\CARRYB[4][9] ), .B(\ab[5][9] ), .ZN(net86102) );
  NAND2_X1 U370 ( .A1(\CARRYB[4][9] ), .A2(\ab[5][9] ), .ZN(net83056) );
  NAND2_X1 U371 ( .A1(\SUMB[4][10] ), .A2(\CARRYB[4][9] ), .ZN(net83054) );
  XNOR2_X1 U372 ( .A(net86070), .B(\SUMB[2][11] ), .ZN(\SUMB[3][10] ) );
  INV_X1 U374 ( .A(A[4]), .ZN(n108) );
  NAND2_X1 U378 ( .A1(net76827), .A2(net76831), .ZN(net110254) );
  CLKBUF_X1 U379 ( .A(ZA), .Z(net76827) );
  CLKBUF_X1 U381 ( .A(net83140), .Z(net77238) );
  NAND2_X1 U382 ( .A1(net83140), .A2(net88254), .ZN(net86087) );
  INV_X1 U384 ( .A(n111), .ZN(n109) );
  CLKBUF_X1 U385 ( .A(TC), .Z(n111) );
  INV_X1 U386 ( .A(A[15]), .ZN(n110) );
  INV_X1 U388 ( .A(B[8]), .ZN(net99186) );
  XNOR2_X1 U391 ( .A(\CARRYB[12][7] ), .B(n112), .ZN(n126) );
  XNOR2_X1 U393 ( .A(n113), .B(\SUMB[15][6] ), .ZN(n36) );
  INV_X1 U395 ( .A(B[11]), .ZN(net94632) );
  NOR2_X1 U397 ( .A1(net94632), .A2(net83231), .ZN(net88235) );
  INV_X1 U399 ( .A(A[2]), .ZN(net97393) );
  INV_X1 U401 ( .A(B[12]), .ZN(net74496) );
  XOR2_X1 U403 ( .A(net83610), .B(net95160), .Z(n21) );
  INV_X1 U404 ( .A(B[12]), .ZN(net82807) );
  CLKBUF_X1 U405 ( .A(A[2]), .Z(net94668) );
  XOR2_X1 U406 ( .A(\CARRYB[14][6] ), .B(\ab[15][6] ), .Z(n114) );
  XOR2_X1 U407 ( .A(\SUMB[14][7] ), .B(n114), .Z(\SUMB[15][6] ) );
  NAND2_X1 U408 ( .A1(\SUMB[14][7] ), .A2(\CARRYB[14][6] ), .ZN(n115) );
  NAND2_X1 U409 ( .A1(\SUMB[14][7] ), .A2(\ab[15][6] ), .ZN(n116) );
  NAND2_X1 U410 ( .A1(\CARRYB[14][6] ), .A2(\ab[15][6] ), .ZN(n117) );
  XNOR2_X1 U413 ( .A(n118), .B(\SUMB[11][6] ), .ZN(\SUMB[12][5] ) );
  XNOR2_X1 U414 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .ZN(n118) );
  CLKBUF_X1 U416 ( .A(net77238), .Z(net112156) );
  XNOR2_X1 U417 ( .A(\SUMB[7][10] ), .B(n119), .ZN(\SUMB[8][9] ) );
  XNOR2_X1 U418 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .ZN(n119) );
  XOR2_X1 U419 ( .A(\ab[4][14] ), .B(\ab[3][15] ), .Z(n120) );
  XOR2_X1 U420 ( .A(\CARRYB[3][14] ), .B(n120), .Z(\SUMB[4][14] ) );
  NAND2_X1 U421 ( .A1(\CARRYB[3][14] ), .A2(\ab[4][14] ), .ZN(n121) );
  NAND2_X1 U422 ( .A1(\CARRYB[3][14] ), .A2(\ab[3][15] ), .ZN(n122) );
  NAND2_X1 U423 ( .A1(\ab[4][14] ), .A2(\ab[3][15] ), .ZN(n123) );
  XNOR2_X1 U426 ( .A(\CARRYB[2][14] ), .B(n125), .ZN(\SUMB[3][14] ) );
  XNOR2_X1 U427 ( .A(\ab[3][14] ), .B(\ab[2][15] ), .ZN(n125) );
  XOR2_X1 U428 ( .A(\SUMB[12][8] ), .B(n126), .Z(\SUMB[13][7] ) );
  NAND2_X1 U429 ( .A1(\SUMB[12][8] ), .A2(\CARRYB[12][7] ), .ZN(n127) );
  NAND2_X1 U430 ( .A1(\SUMB[12][8] ), .A2(\ab[13][7] ), .ZN(n128) );
  NAND2_X1 U431 ( .A1(\CARRYB[12][7] ), .A2(\ab[13][7] ), .ZN(n129) );
  INV_X2 U435 ( .A(B[1]), .ZN(n132) );
  XNOR2_X1 U438 ( .A(net110260), .B(\SUMB[15][1] ), .ZN(n41) );
  XNOR2_X1 U440 ( .A(\SUMB[7][8] ), .B(n134), .ZN(\SUMB[8][7] ) );
  XNOR2_X1 U441 ( .A(\CARRYB[7][7] ), .B(\ab[8][7] ), .ZN(n134) );
  XOR2_X1 U442 ( .A(net76827), .B(net76831), .Z(n135) );
  XOR2_X1 U443 ( .A(\SUMB[15][0] ), .B(n135), .Z(\A1[13] ) );
  XNOR2_X1 U444 ( .A(\SUMB[14][4] ), .B(n136), .ZN(\SUMB[15][3] ) );
  XNOR2_X1 U445 ( .A(\CARRYB[14][3] ), .B(\ab[15][3] ), .ZN(n136) );
  NAND2_X1 U446 ( .A1(\SUMB[14][4] ), .A2(\CARRYB[14][3] ), .ZN(n137) );
  NAND2_X1 U447 ( .A1(\SUMB[14][4] ), .A2(\ab[15][3] ), .ZN(n138) );
  NAND2_X1 U448 ( .A1(\CARRYB[14][3] ), .A2(\ab[15][3] ), .ZN(n139) );
  INV_X1 U450 ( .A(\CARRYB[15][3] ), .ZN(n151) );
  XOR2_X1 U454 ( .A(\CARRYB[13][3] ), .B(\ab[14][3] ), .Z(n140) );
  XOR2_X1 U455 ( .A(n140), .B(\SUMB[13][4] ), .Z(\SUMB[14][3] ) );
  XOR2_X1 U456 ( .A(\CARRYB[14][2] ), .B(\ab[15][2] ), .Z(n141) );
  XOR2_X1 U457 ( .A(n141), .B(\SUMB[14][3] ), .Z(\SUMB[15][2] ) );
  NAND2_X1 U458 ( .A1(\CARRYB[13][3] ), .A2(\ab[14][3] ), .ZN(n142) );
  NAND2_X1 U459 ( .A1(\CARRYB[13][3] ), .A2(\SUMB[13][4] ), .ZN(n143) );
  NAND2_X1 U460 ( .A1(\ab[14][3] ), .A2(\SUMB[13][4] ), .ZN(n144) );
  NAND2_X1 U462 ( .A1(\CARRYB[14][2] ), .A2(\ab[15][2] ), .ZN(n145) );
  NAND2_X1 U463 ( .A1(\CARRYB[14][2] ), .A2(\SUMB[14][3] ), .ZN(n146) );
  NAND2_X1 U464 ( .A1(\ab[15][2] ), .A2(\SUMB[14][3] ), .ZN(n147) );
  CLKBUF_X1 U466 ( .A(net83048), .Z(net95229) );
  XNOR2_X1 U468 ( .A(\SUMB[12][4] ), .B(n148), .ZN(\SUMB[13][3] ) );
  XNOR2_X1 U469 ( .A(\CARRYB[12][3] ), .B(\ab[13][3] ), .ZN(n148) );
  XNOR2_X1 U470 ( .A(n149), .B(n28), .ZN(\SUMB[2][5] ) );
  XNOR2_X1 U471 ( .A(n15), .B(\ab[2][5] ), .ZN(n149) );
  XNOR2_X1 U472 ( .A(n151), .B(\SUMB[15][4] ), .ZN(n150) );
  NAND2_X1 U473 ( .A1(\SUMB[7][10] ), .A2(\CARRYB[7][9] ), .ZN(n152) );
  NAND2_X1 U474 ( .A1(\SUMB[7][10] ), .A2(\ab[8][9] ), .ZN(n153) );
  NAND2_X1 U475 ( .A1(n326), .A2(\ab[8][9] ), .ZN(n154) );
  NAND2_X1 U477 ( .A1(n28), .A2(n15), .ZN(n155) );
  NAND2_X1 U478 ( .A1(n28), .A2(\ab[2][5] ), .ZN(n156) );
  NAND2_X1 U479 ( .A1(n15), .A2(\ab[2][5] ), .ZN(n157) );
  XOR2_X1 U481 ( .A(\CARRYB[10][5] ), .B(\ab[11][5] ), .Z(n158) );
  XOR2_X1 U482 ( .A(\SUMB[10][6] ), .B(n158), .Z(\SUMB[11][5] ) );
  NAND2_X1 U483 ( .A1(\SUMB[10][6] ), .A2(\CARRYB[10][5] ), .ZN(n159) );
  NAND2_X1 U484 ( .A1(\SUMB[10][6] ), .A2(\ab[11][5] ), .ZN(n160) );
  NAND2_X1 U485 ( .A1(\CARRYB[10][5] ), .A2(\ab[11][5] ), .ZN(n161) );
  XNOR2_X1 U487 ( .A(n162), .B(\SUMB[15][3] ), .ZN(n49) );
  XOR2_X1 U489 ( .A(\CARRYB[11][4] ), .B(\ab[12][4] ), .Z(n163) );
  XOR2_X1 U490 ( .A(\SUMB[11][5] ), .B(n163), .Z(\SUMB[12][4] ) );
  NAND2_X1 U491 ( .A1(\SUMB[11][5] ), .A2(\CARRYB[11][4] ), .ZN(n164) );
  NAND2_X1 U492 ( .A1(\SUMB[11][5] ), .A2(\ab[12][4] ), .ZN(n165) );
  NAND2_X1 U493 ( .A1(\CARRYB[11][4] ), .A2(\ab[12][4] ), .ZN(n166) );
  INV_X1 U495 ( .A(net83034), .ZN(net83036) );
  INV_X1 U496 ( .A(B[8]), .ZN(net83624) );
  XOR2_X1 U497 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n30) );
  NAND2_X1 U498 ( .A1(\SUMB[12][4] ), .A2(\CARRYB[12][3] ), .ZN(n167) );
  NAND2_X1 U499 ( .A1(\SUMB[12][4] ), .A2(\ab[13][3] ), .ZN(n168) );
  NAND2_X1 U500 ( .A1(\CARRYB[12][3] ), .A2(\ab[13][3] ), .ZN(n169) );
  XOR2_X1 U502 ( .A(\CARRYB[13][6] ), .B(\ab[14][6] ), .Z(n170) );
  XOR2_X1 U503 ( .A(\SUMB[13][7] ), .B(n170), .Z(\SUMB[14][6] ) );
  NAND2_X1 U504 ( .A1(\SUMB[13][7] ), .A2(\CARRYB[13][6] ), .ZN(n171) );
  NAND2_X1 U505 ( .A1(\SUMB[13][7] ), .A2(\ab[14][6] ), .ZN(n172) );
  NAND2_X1 U506 ( .A1(\CARRYB[13][6] ), .A2(\ab[14][6] ), .ZN(n173) );
  XNOR2_X1 U508 ( .A(\SUMB[6][9] ), .B(n174), .ZN(\SUMB[7][8] ) );
  XNOR2_X1 U509 ( .A(\CARRYB[6][8] ), .B(\ab[7][8] ), .ZN(n174) );
  XNOR2_X1 U513 ( .A(n176), .B(n25), .ZN(\SUMB[2][11] ) );
  XNOR2_X1 U514 ( .A(\ab[2][11] ), .B(n9), .ZN(n176) );
  XNOR2_X1 U515 ( .A(\SUMB[10][9] ), .B(n177), .ZN(\SUMB[11][8] ) );
  XNOR2_X1 U516 ( .A(\CARRYB[10][8] ), .B(\ab[11][8] ), .ZN(n177) );
  XNOR2_X1 U518 ( .A(\SUMB[15][5] ), .B(n179), .ZN(n50) );
  INV_X1 U520 ( .A(B[13]), .ZN(net86104) );
  XNOR2_X1 U521 ( .A(net86102), .B(\SUMB[4][10] ), .ZN(\SUMB[5][9] ) );
  NAND2_X1 U522 ( .A1(net88201), .A2(n183), .ZN(n180) );
  NAND2_X1 U523 ( .A1(n180), .A2(n181), .ZN(n17) );
  OR2_X1 U524 ( .A1(n205), .A2(net86087), .ZN(n181) );
  NAND2_X1 U527 ( .A1(\SUMB[6][9] ), .A2(\CARRYB[6][8] ), .ZN(n184) );
  NAND2_X1 U528 ( .A1(\SUMB[6][9] ), .A2(\ab[7][8] ), .ZN(n185) );
  NAND2_X1 U529 ( .A1(\CARRYB[6][8] ), .A2(\ab[7][8] ), .ZN(n186) );
  NAND2_X1 U531 ( .A1(\SUMB[10][9] ), .A2(\CARRYB[10][8] ), .ZN(n187) );
  NAND2_X1 U532 ( .A1(\SUMB[10][9] ), .A2(\ab[11][8] ), .ZN(n188) );
  NAND2_X1 U533 ( .A1(\CARRYB[10][8] ), .A2(\ab[11][8] ), .ZN(n189) );
  NAND2_X1 U535 ( .A1(\SUMB[7][8] ), .A2(\CARRYB[7][7] ), .ZN(n190) );
  NAND2_X1 U536 ( .A1(\SUMB[7][8] ), .A2(\ab[8][7] ), .ZN(n191) );
  NAND2_X1 U537 ( .A1(\CARRYB[7][7] ), .A2(\ab[8][7] ), .ZN(n192) );
  INV_X1 U540 ( .A(n193), .ZN(n205) );
  NAND2_X1 U541 ( .A1(\ab[2][11] ), .A2(n9), .ZN(n194) );
  NAND2_X1 U542 ( .A1(\ab[2][11] ), .A2(n25), .ZN(n195) );
  NAND2_X1 U543 ( .A1(n9), .A2(n25), .ZN(n196) );
  NAND2_X1 U545 ( .A1(\CARRYB[2][10] ), .A2(\ab[3][10] ), .ZN(n197) );
  NAND2_X1 U546 ( .A1(\SUMB[2][11] ), .A2(\CARRYB[2][10] ), .ZN(n198) );
  NAND2_X1 U547 ( .A1(\SUMB[2][11] ), .A2(\ab[3][10] ), .ZN(n199) );
  XNOR2_X1 U553 ( .A(n200), .B(\SUMB[8][10] ), .ZN(\SUMB[9][9] ) );
  XNOR2_X1 U554 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .ZN(n200) );
  INV_X1 U559 ( .A(B[5]), .ZN(n318) );
  INV_X1 U560 ( .A(B[11]), .ZN(net82848) );
  INV_X1 U562 ( .A(\SUMB[2][4] ), .ZN(n209) );
  XNOR2_X1 U564 ( .A(n204), .B(\ab[0][14] ), .ZN(n26) );
  OR2_X1 U565 ( .A1(net86104), .A2(net83231), .ZN(n204) );
  INV_X1 U571 ( .A(B[14]), .ZN(net83506) );
  NOR2_X1 U574 ( .A1(net86104), .A2(net83230), .ZN(n207) );
  XNOR2_X1 U577 ( .A(n209), .B(n245), .ZN(\SUMB[3][3] ) );
  INV_X1 U578 ( .A(net82807), .ZN(net83413) );
  INV_X2 U580 ( .A(net83413), .ZN(net83415) );
  CLKBUF_X1 U581 ( .A(net74499), .Z(net83407) );
  XNOR2_X1 U582 ( .A(n210), .B(\SUMB[7][11] ), .ZN(\SUMB[8][10] ) );
  XNOR2_X1 U583 ( .A(\CARRYB[7][10] ), .B(\ab[8][10] ), .ZN(n210) );
  XNOR2_X1 U585 ( .A(\SUMB[10][7] ), .B(n211), .ZN(\SUMB[11][6] ) );
  XNOR2_X1 U586 ( .A(\CARRYB[10][6] ), .B(\ab[11][6] ), .ZN(n211) );
  NAND2_X1 U587 ( .A1(B[7]), .A2(net88197), .ZN(net83284) );
  XNOR2_X1 U588 ( .A(n212), .B(n220), .ZN(\SUMB[4][12] ) );
  INV_X1 U589 ( .A(\SUMB[3][13] ), .ZN(n212) );
  NAND2_X1 U590 ( .A1(\ab[8][10] ), .A2(\CARRYB[7][10] ), .ZN(n213) );
  NAND2_X1 U591 ( .A1(\SUMB[7][11] ), .A2(\ab[8][10] ), .ZN(n214) );
  NAND2_X1 U592 ( .A1(\SUMB[7][11] ), .A2(\CARRYB[7][10] ), .ZN(n215) );
  NAND2_X1 U594 ( .A1(\ab[9][9] ), .A2(\CARRYB[8][9] ), .ZN(n216) );
  NAND2_X1 U595 ( .A1(n327), .A2(\ab[9][9] ), .ZN(n217) );
  NAND2_X1 U596 ( .A1(n327), .A2(\CARRYB[8][9] ), .ZN(n218) );
  XNOR2_X1 U598 ( .A(\CARRYB[2][3] ), .B(n219), .ZN(n245) );
  INV_X1 U600 ( .A(A[1]), .ZN(net83230) );
  XOR2_X1 U603 ( .A(\CARRYB[3][12] ), .B(\ab[4][12] ), .Z(n220) );
  NAND2_X1 U604 ( .A1(\SUMB[3][13] ), .A2(\CARRYB[3][12] ), .ZN(n221) );
  NAND2_X1 U605 ( .A1(\SUMB[3][13] ), .A2(\ab[4][12] ), .ZN(n222) );
  NAND2_X1 U606 ( .A1(\CARRYB[3][12] ), .A2(\ab[4][12] ), .ZN(n223) );
  XNOR2_X1 U608 ( .A(\ab[0][15] ), .B(n205), .ZN(n224) );
  XNOR2_X1 U609 ( .A(n224), .B(n260), .ZN(n225) );
  XNOR2_X1 U610 ( .A(\SUMB[6][11] ), .B(n226), .ZN(\SUMB[7][10] ) );
  CLKBUF_X1 U612 ( .A(net86104), .Z(net83154) );
  XOR2_X1 U615 ( .A(\CARRYB[5][10] ), .B(\ab[6][10] ), .Z(n228) );
  XOR2_X1 U616 ( .A(n228), .B(\SUMB[5][11] ), .Z(\SUMB[6][10] ) );
  NAND2_X1 U617 ( .A1(\SUMB[5][11] ), .A2(n325), .ZN(n229) );
  NAND2_X1 U618 ( .A1(\SUMB[5][11] ), .A2(\ab[6][10] ), .ZN(n230) );
  NAND2_X1 U619 ( .A1(n325), .A2(\ab[6][10] ), .ZN(n231) );
  XNOR2_X1 U623 ( .A(\SUMB[9][6] ), .B(net83091), .ZN(\SUMB[10][5] ) );
  XNOR2_X1 U624 ( .A(\SUMB[5][9] ), .B(net83077), .ZN(\SUMB[6][8] ) );
  XNOR2_X1 U625 ( .A(\ab[0][15] ), .B(n205), .ZN(n31) );
  NAND2_X1 U626 ( .A1(\SUMB[4][10] ), .A2(\ab[5][9] ), .ZN(n233) );
  NAND2_X1 U628 ( .A1(\SUMB[9][6] ), .A2(\ab[10][5] ), .ZN(n234) );
  NAND2_X1 U630 ( .A1(\SUMB[10][7] ), .A2(\CARRYB[10][6] ), .ZN(n235) );
  NAND2_X1 U631 ( .A1(\SUMB[10][7] ), .A2(\ab[11][6] ), .ZN(n236) );
  NAND2_X1 U632 ( .A1(\CARRYB[10][6] ), .A2(\ab[11][6] ), .ZN(n237) );
  XNOR2_X1 U635 ( .A(n239), .B(\SUMB[4][12] ), .ZN(\SUMB[5][11] ) );
  XNOR2_X1 U636 ( .A(\CARRYB[4][11] ), .B(\ab[5][11] ), .ZN(n239) );
  XOR2_X1 U637 ( .A(\SUMB[13][1] ), .B(\ab[14][0] ), .Z(n240) );
  XOR2_X1 U638 ( .A(\CARRYB[13][0] ), .B(n240), .Z(\A1[12] ) );
  NAND2_X1 U639 ( .A1(\CARRYB[13][0] ), .A2(\SUMB[13][1] ), .ZN(n241) );
  NAND2_X1 U640 ( .A1(\CARRYB[13][0] ), .A2(\ab[14][0] ), .ZN(n242) );
  NAND2_X1 U641 ( .A1(\SUMB[13][1] ), .A2(\ab[14][0] ), .ZN(n243) );
  NAND2_X1 U644 ( .A1(\SUMB[5][9] ), .A2(\ab[6][8] ), .ZN(n244) );
  NAND2_X1 U646 ( .A1(\SUMB[2][4] ), .A2(\CARRYB[2][3] ), .ZN(n246) );
  NAND2_X1 U647 ( .A1(\SUMB[2][4] ), .A2(\ab[3][3] ), .ZN(n247) );
  NAND2_X1 U648 ( .A1(\CARRYB[2][3] ), .A2(\ab[3][3] ), .ZN(n248) );
  XNOR2_X1 U650 ( .A(net83153), .B(n249), .ZN(n25) );
  OR2_X1 U651 ( .A1(net82807), .A2(net83231), .ZN(n249) );
  XNOR2_X1 U652 ( .A(n250), .B(\SUMB[6][10] ), .ZN(\SUMB[7][9] ) );
  XNOR2_X1 U653 ( .A(\CARRYB[6][9] ), .B(\ab[7][9] ), .ZN(n250) );
  NAND2_X1 U654 ( .A1(\SUMB[11][6] ), .A2(\CARRYB[11][5] ), .ZN(n251) );
  NAND2_X1 U655 ( .A1(\SUMB[11][6] ), .A2(\ab[12][5] ), .ZN(n252) );
  NAND2_X1 U656 ( .A1(\CARRYB[11][5] ), .A2(\ab[12][5] ), .ZN(n253) );
  NAND2_X1 U658 ( .A1(\SUMB[6][11] ), .A2(n324), .ZN(n254) );
  NAND2_X1 U659 ( .A1(\SUMB[6][11] ), .A2(\ab[7][10] ), .ZN(n255) );
  NAND2_X1 U660 ( .A1(n324), .A2(\ab[7][10] ), .ZN(n256) );
  NAND2_X1 U662 ( .A1(\CARRYB[2][14] ), .A2(\ab[3][14] ), .ZN(n257) );
  NAND2_X1 U663 ( .A1(\CARRYB[2][14] ), .A2(\ab[2][15] ), .ZN(n258) );
  NAND2_X1 U664 ( .A1(\ab[3][14] ), .A2(\ab[2][15] ), .ZN(n259) );
  XNOR2_X1 U666 ( .A(n224), .B(n260), .ZN(\SUMB[2][13] ) );
  XNOR2_X1 U667 ( .A(\ab[2][13] ), .B(n12), .ZN(n260) );
  NOR2_X1 U668 ( .A1(net74499), .A2(TC), .ZN(net82786) );
  NOR2_X1 U669 ( .A1(net83231), .A2(net82807), .ZN(n261) );
  INV_X1 U670 ( .A(net83407), .ZN(net82665) );
  XNOR2_X1 U671 ( .A(n262), .B(\SUMB[2][13] ), .ZN(\SUMB[3][12] ) );
  XNOR2_X1 U672 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .ZN(n262) );
  NAND2_X1 U673 ( .A1(n31), .A2(\ab[2][13] ), .ZN(n263) );
  NAND2_X1 U674 ( .A1(n31), .A2(n12), .ZN(n264) );
  NAND2_X1 U675 ( .A1(\ab[2][13] ), .A2(n12), .ZN(n265) );
  NAND2_X1 U677 ( .A1(\SUMB[4][12] ), .A2(\CARRYB[4][11] ), .ZN(n266) );
  NAND2_X1 U678 ( .A1(\SUMB[4][12] ), .A2(\ab[5][11] ), .ZN(n267) );
  NAND2_X1 U679 ( .A1(\CARRYB[4][11] ), .A2(\ab[5][11] ), .ZN(n268) );
  NAND2_X1 U681 ( .A1(\CARRYB[6][9] ), .A2(\SUMB[6][10] ), .ZN(n269) );
  NAND2_X1 U682 ( .A1(\SUMB[6][10] ), .A2(\ab[7][9] ), .ZN(n270) );
  NAND2_X1 U683 ( .A1(\CARRYB[6][9] ), .A2(\ab[7][9] ), .ZN(n271) );
  NAND2_X1 U685 ( .A1(\SUMB[6][8] ), .A2(\CARRYB[6][7] ), .ZN(n272) );
  NAND2_X1 U686 ( .A1(\SUMB[6][8] ), .A2(\ab[7][7] ), .ZN(n273) );
  INV_X1 U688 ( .A(\CARRYB[15][1] ), .ZN(net82656) );
  XNOR2_X1 U689 ( .A(\SUMB[15][2] ), .B(net82656), .ZN(n34) );
  NAND2_X1 U690 ( .A1(\SUMB[11][4] ), .A2(\ab[12][3] ), .ZN(n274) );
  NAND2_X1 U692 ( .A1(\SUMB[2][13] ), .A2(\CARRYB[2][12] ), .ZN(n275) );
  NAND2_X1 U693 ( .A1(n225), .A2(\ab[3][12] ), .ZN(n276) );
  NAND2_X1 U694 ( .A1(\CARRYB[2][12] ), .A2(\ab[3][12] ), .ZN(n277) );
  CLKBUF_X1 U696 ( .A(n319), .Z(n303) );
  CLKBUF_X1 U697 ( .A(n320), .Z(n306) );
  INV_X1 U728 ( .A(B[4]), .ZN(n319) );
  INV_X1 U729 ( .A(B[3]), .ZN(n320) );
  INV_X1 U730 ( .A(A[7]), .ZN(n315) );
  INV_X1 U731 ( .A(A[11]), .ZN(n312) );
  INV_X1 U732 ( .A(A[14]), .ZN(n310) );
  INV_X1 U733 ( .A(A[6]), .ZN(n316) );
  INV_X1 U734 ( .A(A[10]), .ZN(n313) );
  INV_X1 U735 ( .A(A[12]), .ZN(n311) );
  INV_X1 U736 ( .A(A[5]), .ZN(n317) );
  INV_X1 U737 ( .A(A[9]), .ZN(n314) );
  INV_X1 U738 ( .A(B[0]), .ZN(n322) );
  INV_X1 U739 ( .A(B[15]), .ZN(net74499) );
  ALU_N32_DW01_add_0 FS_1 ( .A({n63, n62, n40, n54, n39, n53, n38, n52, n37, 
        n51, n36, n50, n150, n49, n34, n41, \A1[13] , \A1[12] , \A1[11] , 
        \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , 
        \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n32, n61, n48, n60, n47, n59, 
        n46, n58, n45, n57, n44, n56, n43, n55, n42, \A2[14] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[31:2]) );
  AND2_X1 U2 ( .A1(\ab[0][12] ), .A2(net88235), .ZN(n9) );
  BUF_X1 U3 ( .A(n108), .Z(net76873) );
  BUF_X1 U4 ( .A(n108), .Z(net76872) );
  BUF_X1 U5 ( .A(net82786), .Z(net76821) );
  INV_X1 U7 ( .A(net94668), .ZN(net83786) );
  AND2_X1 U8 ( .A1(\SUMB[15][1] ), .A2(\CARRYB[15][0] ), .ZN(n42) );
  AND2_X1 U9 ( .A1(\CARRYB[15][4] ), .A2(\SUMB[15][5] ), .ZN(n44) );
  MUX2_X1 U10 ( .A(net76821), .B(net76831), .S(net83786), .Z(\ab[2][15] ) );
  MUX2_X2 U11 ( .A(net82786), .B(net83140), .S(net82901), .Z(\ab[0][15] ) );
  AND2_X1 U12 ( .A1(B[2]), .A2(net88197), .ZN(n323) );
  AND2_X1 U13 ( .A1(B[15]), .A2(TC), .ZN(net83140) );
  CLKBUF_X1 U14 ( .A(\CARRYB[6][10] ), .Z(n324) );
  BUF_X1 U15 ( .A(\CARRYB[5][10] ), .Z(n325) );
  NAND3_X1 U16 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n326) );
  XNOR2_X1 U20 ( .A(n210), .B(\SUMB[7][11] ), .ZN(n327) );
  XNOR2_X1 U22 ( .A(\CARRYB[6][10] ), .B(\ab[7][10] ), .ZN(n226) );
  BUF_X2 U23 ( .A(net83140), .Z(net76831) );
  XOR2_X1 U29 ( .A(\CARRYB[2][13] ), .B(\ab[3][13] ), .Z(n328) );
  XOR2_X1 U31 ( .A(\SUMB[2][14] ), .B(n328), .Z(\SUMB[3][13] ) );
  NAND2_X1 U33 ( .A1(\SUMB[2][14] ), .A2(\CARRYB[2][13] ), .ZN(n329) );
  NAND2_X1 U35 ( .A1(\SUMB[2][14] ), .A2(\ab[3][13] ), .ZN(n330) );
  NAND2_X1 U43 ( .A1(\CARRYB[2][13] ), .A2(\ab[3][13] ), .ZN(n331) );
  NAND3_X1 U44 ( .A1(n329), .A2(n330), .A3(n331), .ZN(\CARRYB[3][13] ) );
  BUF_X1 U45 ( .A(net74503), .Z(net76865) );
  MUX2_X1 U46 ( .A(net76821), .B(net76831), .S(n315), .Z(\ab[7][15] ) );
  AND2_X1 U47 ( .A1(\CARRYB[15][9] ), .A2(\SUMB[15][10] ), .ZN(n59) );
  CLKBUF_X1 U48 ( .A(net82786), .Z(net88201) );
  NAND3_X1 U49 ( .A1(n263), .A2(n264), .A3(n265), .ZN(\CARRYB[2][13] ) );
  NAND3_X1 U56 ( .A1(n194), .A2(n195), .A3(n196), .ZN(\CARRYB[2][11] ) );
  MUX2_X1 U57 ( .A(net76821), .B(net76831), .S(net76872), .Z(\ab[4][15] ) );
  NAND3_X1 U58 ( .A1(n121), .A2(n122), .A3(n123), .ZN(\CARRYB[4][14] ) );
  NAND3_X1 U59 ( .A1(net83054), .A2(n233), .A3(net83056), .ZN(\CARRYB[5][9] )
         );
  NAND3_X1 U60 ( .A1(n214), .A2(n213), .A3(n215), .ZN(\CARRYB[8][10] ) );
  MUX2_X1 U61 ( .A(net76821), .B(net76831), .S(n314), .Z(\ab[9][15] ) );
  NAND3_X1 U62 ( .A1(n142), .A2(n143), .A3(n144), .ZN(\CARRYB[14][3] ) );
  NAND3_X1 U67 ( .A1(n187), .A2(n188), .A3(n189), .ZN(\CARRYB[11][8] ) );
  NAND3_X1 U68 ( .A1(n235), .A2(n236), .A3(n237), .ZN(\CARRYB[11][6] ) );
  MUX2_X1 U69 ( .A(net76821), .B(net112156), .S(n311), .Z(\ab[12][15] ) );
  MUX2_X1 U70 ( .A(n99), .B(ZA), .S(n132), .Z(\ab[15][1] ) );
  MUX2_X1 U71 ( .A(n99), .B(net76827), .S(net83036), .Z(\ab[15][9] ) );
  MUX2_X1 U72 ( .A(n99), .B(ZA), .S(net95229), .Z(\ab[15][10] ) );
  AND2_X1 U75 ( .A1(\CARRYB[15][11] ), .A2(\SUMB[15][12] ), .ZN(n60) );
  AND2_X1 U78 ( .A1(B[14]), .A2(net88197), .ZN(n193) );
  AND2_X1 U80 ( .A1(B[14]), .A2(net82934), .ZN(\ab[0][14] ) );
  MUX2_X1 U81 ( .A(net88201), .B(net77238), .S(net83230), .Z(\ab[1][15] ) );
  AND2_X1 U82 ( .A1(A[1]), .A2(B[10]), .ZN(net95160) );
  NAND3_X1 U87 ( .A1(n275), .A2(n276), .A3(n277), .ZN(\CARRYB[3][12] ) );
  MUX2_X1 U88 ( .A(net76821), .B(net76831), .S(n316), .Z(\ab[6][15] ) );
  AND2_X1 U92 ( .A1(B[8]), .A2(net88197), .ZN(\ab[1][8] ) );
  NAND3_X1 U95 ( .A1(n229), .A2(n230), .A3(n231), .ZN(\CARRYB[6][10] ) );
  NAND3_X1 U96 ( .A1(n266), .A2(n267), .A3(n268), .ZN(\CARRYB[5][11] ) );
  NAND3_X1 U107 ( .A1(n272), .A2(n273), .A3(net82664), .ZN(\CARRYB[7][7] ) );
  NAND3_X1 U123 ( .A1(n184), .A2(n185), .A3(n186), .ZN(\CARRYB[7][8] ) );
  AND2_X1 U139 ( .A1(\ab[1][6] ), .A2(\ab[0][7] ), .ZN(n14) );
  AND2_X1 U155 ( .A1(B[6]), .A2(net94668), .ZN(\ab[2][6] ) );
  NAND3_X1 U171 ( .A1(net83042), .A2(n234), .A3(net83044), .ZN(\CARRYB[10][5] ) );
  NAND3_X1 U187 ( .A1(n152), .A2(n153), .A3(n154), .ZN(\CARRYB[8][9] ) );
  AND2_X1 U203 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n15) );
  NAND3_X1 U213 ( .A1(n167), .A2(n168), .A3(n169), .ZN(\CARRYB[13][3] ) );
  MUX2_X1 U219 ( .A(net76821), .B(net112156), .S(n313), .Z(\ab[10][15] ) );
  MUX2_X1 U228 ( .A(n99), .B(ZA), .S(net74486), .Z(\ab[15][2] ) );
  MUX2_X1 U235 ( .A(n99), .B(ZA), .S(n320), .Z(\ab[15][3] ) );
  NAND3_X1 U237 ( .A1(n164), .A2(n165), .A3(n166), .ZN(\CARRYB[12][4] ) );
  NAND3_X1 U238 ( .A1(n251), .A2(n252), .A3(n253), .ZN(\CARRYB[12][5] ) );
  AND2_X1 U239 ( .A1(\ab[1][3] ), .A2(\ab[0][4] ), .ZN(n3) );
  AND2_X1 U240 ( .A1(\ab[1][4] ), .A2(\ab[0][5] ), .ZN(n16) );
  INV_X1 U242 ( .A(B[5]), .ZN(n201) );
  INV_X1 U243 ( .A(\ab[13][7] ), .ZN(n112) );
  NAND3_X1 U244 ( .A1(net110252), .A2(net110253), .A3(net110254), .ZN(\A2[14] ) );
  INV_X1 U245 ( .A(\CARRYB[15][0] ), .ZN(net110260) );
  INV_X1 U246 ( .A(\CARRYB[15][2] ), .ZN(n162) );
  AND2_X1 U247 ( .A1(\CARRYB[15][1] ), .A2(\SUMB[15][2] ), .ZN(n55) );
  INV_X1 U248 ( .A(\CARRYB[15][4] ), .ZN(n179) );
  AND2_X1 U249 ( .A1(\CARRYB[15][3] ), .A2(\SUMB[15][4] ), .ZN(n56) );
  INV_X1 U250 ( .A(\CARRYB[15][5] ), .ZN(n113) );
  NAND3_X1 U252 ( .A1(n115), .A2(n116), .A3(n117), .ZN(\CARRYB[15][6] ) );
  MUX2_X1 U253 ( .A(n99), .B(net76827), .S(net83313), .Z(\ab[15][7] ) );
  AND2_X1 U254 ( .A1(\SUMB[15][6] ), .A2(\CARRYB[15][5] ), .ZN(n57) );
  MUX2_X1 U255 ( .A(net76821), .B(net76831), .S(n102), .Z(\ab[13][15] ) );
  AND2_X1 U256 ( .A1(\CARRYB[15][6] ), .A2(\SUMB[15][7] ), .ZN(n45) );
  MUX2_X1 U257 ( .A(n99), .B(ZA), .S(net82848), .Z(\ab[15][11] ) );
  AND2_X1 U268 ( .A1(\CARRYB[15][13] ), .A2(\SUMB[15][14] ), .ZN(n61) );
  MUX2_X1 U284 ( .A(n99), .B(ZA), .S(net83415), .Z(\ab[15][12] ) );
  AND2_X1 U300 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n4) );
  AND2_X1 U316 ( .A1(\CARRYB[15][10] ), .A2(\SUMB[15][11] ), .ZN(n47) );
  AND2_X1 U332 ( .A1(n207), .A2(\ab[0][14] ), .ZN(n12) );
  AND2_X1 U341 ( .A1(net82934), .A2(n193), .ZN(n183) );
  AND2_X1 U348 ( .A1(net83153), .A2(n261), .ZN(n11) );
  NAND3_X1 U351 ( .A1(n257), .A2(n258), .A3(n259), .ZN(\CARRYB[3][14] ) );
  MUX2_X1 U353 ( .A(net76821), .B(net77238), .S(net76866), .Z(\ab[3][15] ) );
  MUX2_X1 U359 ( .A(net76821), .B(net76831), .S(n317), .Z(\ab[5][15] ) );
  AND2_X1 U364 ( .A1(net97340), .A2(net83498), .ZN(n10) );
  AND2_X1 U373 ( .A1(net83034), .A2(net94668), .ZN(\ab[2][9] ) );
  NAND3_X1 U375 ( .A1(n197), .A2(n198), .A3(n199), .ZN(\CARRYB[3][10] ) );
  NAND3_X1 U376 ( .A1(n221), .A2(n222), .A3(n223), .ZN(\CARRYB[4][12] ) );
  AND2_X1 U377 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n8) );
  NAND3_X1 U380 ( .A1(net82866), .A2(n244), .A3(net82868), .ZN(\CARRYB[6][8] )
         );
  AND2_X1 U383 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n13) );
  NAND3_X1 U387 ( .A1(n254), .A2(n255), .A3(n256), .ZN(\CARRYB[7][10] ) );
  NAND3_X1 U389 ( .A1(n269), .A2(n270), .A3(n271), .ZN(\CARRYB[7][9] ) );
  MUX2_X1 U390 ( .A(net76821), .B(net76831), .S(net74508), .Z(\ab[8][15] ) );
  AND2_X1 U392 ( .A1(net82934), .A2(B[7]), .ZN(\ab[0][7] ) );
  AND2_X1 U394 ( .A1(B[6]), .A2(net88197), .ZN(\ab[1][6] ) );
  NAND3_X1 U396 ( .A1(n190), .A2(n191), .A3(n192), .ZN(\CARRYB[8][7] ) );
  NAND3_X1 U398 ( .A1(n156), .A2(n155), .A3(n157), .ZN(\CARRYB[2][5] ) );
  NAND3_X1 U400 ( .A1(n160), .A2(n159), .A3(n161), .ZN(\CARRYB[11][5] ) );
  NAND3_X1 U402 ( .A1(n216), .A2(n217), .A3(n218), .ZN(\CARRYB[9][9] ) );
  AND2_X1 U411 ( .A1(B[6]), .A2(net82934), .ZN(\ab[0][6] ) );
  NAND3_X1 U412 ( .A1(net82644), .A2(n274), .A3(net82646), .ZN(\CARRYB[12][3] ) );
  MUX2_X1 U415 ( .A(net76821), .B(net76831), .S(n312), .Z(\ab[11][15] ) );
  BUF_X1 U424 ( .A(A[1]), .Z(net88197) );
  INV_X1 U425 ( .A(\ab[3][3] ), .ZN(n219) );
  NAND3_X1 U432 ( .A1(n246), .A2(n247), .A3(n248), .ZN(\CARRYB[3][3] ) );
  NAND3_X1 U433 ( .A1(n137), .A2(n138), .A3(n139), .ZN(\CARRYB[15][3] ) );
  NAND3_X1 U434 ( .A1(n145), .A2(n146), .A3(n147), .ZN(\CARRYB[15][2] ) );
  NAND3_X1 U436 ( .A1(n171), .A2(n172), .A3(n173), .ZN(\CARRYB[14][6] ) );
  MUX2_X1 U437 ( .A(n99), .B(net76827), .S(net83346), .Z(\ab[15][6] ) );
  NAND3_X1 U439 ( .A1(n127), .A2(n128), .A3(n129), .ZN(\CARRYB[13][7] ) );
  AND2_X1 U449 ( .A1(\CARRYB[15][2] ), .A2(\SUMB[15][3] ), .ZN(n43) );
  MUX2_X1 U451 ( .A(n99), .B(ZA), .S(n303), .Z(\ab[15][4] ) );
  MUX2_X1 U452 ( .A(n99), .B(ZA), .S(n201), .Z(\ab[15][5] ) );
  MUX2_X1 U453 ( .A(n99), .B(net76827), .S(net83624), .Z(\ab[15][8] ) );
  AND2_X1 U461 ( .A1(\CARRYB[15][7] ), .A2(\SUMB[15][8] ), .ZN(n58) );
  BUF_X1 U465 ( .A(net83058), .Z(net88254) );
  AND2_X1 U467 ( .A1(\ab[0][3] ), .A2(n323), .ZN(n5) );
  AND2_X1 U476 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n6) );
  MUX2_X1 U480 ( .A(n99), .B(ZA), .S(n322), .Z(\ab[15][0] ) );
  NAND3_X1 U486 ( .A1(n241), .A2(n243), .A3(n242), .ZN(\CARRYB[14][0] ) );
  AND2_X1 U488 ( .A1(\CARRYB[15][8] ), .A2(\SUMB[15][9] ), .ZN(n46) );
  MUX2_X1 U494 ( .A(net76821), .B(net112156), .S(n310), .Z(\ab[14][15] ) );
  MUX2_X1 U501 ( .A(n99), .B(ZA), .S(net83506), .Z(\ab[15][14] ) );
  MUX2_X1 U507 ( .A(n99), .B(ZA), .S(net83154), .Z(\ab[15][13] ) );
  AND2_X1 U510 ( .A1(\CARRYB[15][14] ), .A2(\SUMB[15][15] ), .ZN(n32) );
  AND2_X1 U511 ( .A1(\CARRYB[15][12] ), .A2(\SUMB[15][13] ), .ZN(n48) );
endmodule


module ALU_N32_DW01_addsub_2 ( A, B, CI, ADD_SUB, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353;

  CLKBUF_X1 U2 ( .A(ADD_SUB), .Z(n353) );
  AND2_X1 U3 ( .A1(n75), .A2(n62), .ZN(n1) );
  AND2_X1 U4 ( .A1(n192), .A2(n193), .ZN(n2) );
  AND2_X1 U5 ( .A1(n277), .A2(n278), .ZN(n3) );
  AND2_X1 U6 ( .A1(n113), .A2(n114), .ZN(n4) );
  AND2_X1 U7 ( .A1(n329), .A2(n45), .ZN(n5) );
  AND2_X1 U8 ( .A1(n114), .A2(n115), .ZN(n6) );
  CLKBUF_X1 U9 ( .A(ADD_SUB), .Z(n352) );
  AOI21_X1 U10 ( .B1(n284), .B2(n12), .A(n285), .ZN(n281) );
  XNOR2_X1 U11 ( .A(B[21]), .B(n352), .ZN(n180) );
  AOI21_X1 U12 ( .B1(n337), .B2(n96), .A(n338), .ZN(n333) );
  AOI21_X1 U13 ( .B1(n316), .B2(n30), .A(n317), .ZN(n312) );
  XNOR2_X1 U14 ( .A(B[9]), .B(n353), .ZN(n301) );
  XNOR2_X1 U15 ( .A(B[11]), .B(n353), .ZN(n294) );
  XNOR2_X1 U16 ( .A(B[12]), .B(n353), .ZN(n287) );
  XNOR2_X1 U17 ( .A(B[13]), .B(n353), .ZN(n272) );
  XNOR2_X1 U18 ( .A(B[14]), .B(n353), .ZN(n265) );
  XNOR2_X1 U19 ( .A(B[15]), .B(n353), .ZN(n257) );
  OAI21_X1 U20 ( .B1(n281), .B2(n282), .A(n283), .ZN(n280) );
  NOR2_X1 U21 ( .A1(n237), .A2(n238), .ZN(n235) );
  NAND4_X1 U22 ( .A1(n12), .A2(n16), .A3(n286), .A4(n279), .ZN(n243) );
  XNOR2_X1 U23 ( .A(B[16]), .B(n352), .ZN(n252) );
  XNOR2_X1 U24 ( .A(B[18]), .B(n352), .ZN(n215) );
  XNOR2_X1 U25 ( .A(B[17]), .B(n352), .ZN(n219) );
  XNOR2_X1 U26 ( .A(B[20]), .B(n352), .ZN(n187) );
  XNOR2_X1 U27 ( .A(B[23]), .B(n352), .ZN(n165) );
  NAND2_X1 U28 ( .A1(A[21]), .A2(n179), .ZN(n177) );
  XNOR2_X1 U29 ( .A(B[22]), .B(n352), .ZN(n173) );
  NAND2_X1 U30 ( .A1(A[24]), .A2(n145), .ZN(n143) );
  NAND2_X1 U31 ( .A1(A[25]), .A2(n138), .ZN(n136) );
  XNOR2_X1 U32 ( .A(B[25]), .B(n352), .ZN(n139) );
  XNOR2_X1 U33 ( .A(B[24]), .B(n352), .ZN(n146) );
  XNOR2_X1 U34 ( .A(B[27]), .B(n352), .ZN(n126) );
  XNOR2_X1 U35 ( .A(B[26]), .B(n352), .ZN(n132) );
  XNOR2_X1 U36 ( .A(B[0]), .B(n353), .ZN(n348) );
  XNOR2_X1 U37 ( .A(B[29]), .B(n352), .ZN(n101) );
  XNOR2_X1 U38 ( .A(B[30]), .B(n352), .ZN(n88) );
  AOI21_X1 U39 ( .B1(n198), .B2(n71), .A(n199), .ZN(n195) );
  NAND2_X1 U40 ( .A1(n187), .A2(n188), .ZN(n161) );
  INV_X1 U41 ( .A(A[20]), .ZN(n188) );
  NAND2_X1 U42 ( .A1(n180), .A2(n181), .ZN(n159) );
  INV_X1 U43 ( .A(A[21]), .ZN(n181) );
  NAND2_X1 U44 ( .A1(A[22]), .A2(n172), .ZN(n157) );
  XNOR2_X1 U45 ( .A(B[19]), .B(n352), .ZN(n209) );
  XNOR2_X1 U46 ( .A(B[1]), .B(n353), .ZN(n340) );
  XNOR2_X1 U47 ( .A(B[2]), .B(n353), .ZN(n335) );
  XNOR2_X1 U48 ( .A(B[3]), .B(n353), .ZN(n331) );
  XNOR2_X1 U49 ( .A(B[4]), .B(n353), .ZN(n321) );
  OAI21_X1 U50 ( .B1(n333), .B2(n41), .A(n42), .ZN(n332) );
  NAND2_X1 U51 ( .A1(n352), .A2(n245), .ZN(n203) );
  XNOR2_X1 U52 ( .A(B[5]), .B(n353), .ZN(n319) );
  XNOR2_X1 U53 ( .A(B[6]), .B(n353), .ZN(n315) );
  XNOR2_X1 U54 ( .A(B[7]), .B(n353), .ZN(n310) );
  XNOR2_X1 U55 ( .A(B[8]), .B(n353), .ZN(n304) );
  NAND2_X1 U56 ( .A1(n308), .A2(n25), .ZN(n251) );
  OAI21_X1 U57 ( .B1(n312), .B2(n313), .A(n21), .ZN(n311) );
  NAND4_X1 U58 ( .A1(n36), .A2(n24), .A3(n30), .A4(n22), .ZN(n242) );
  NAND2_X1 U59 ( .A1(A[9]), .A2(n300), .ZN(n13) );
  NAND2_X1 U60 ( .A1(n301), .A2(n343), .ZN(n12) );
  INV_X1 U61 ( .A(A[9]), .ZN(n343) );
  NAND2_X1 U62 ( .A1(n302), .A2(n17), .ZN(n11) );
  NAND2_X1 U63 ( .A1(n15), .A2(n16), .ZN(n302) );
  XNOR2_X1 U64 ( .A(B[10]), .B(n353), .ZN(n344) );
  NAND2_X1 U65 ( .A1(A[11]), .A2(n296), .ZN(n278) );
  NAND2_X1 U66 ( .A1(n294), .A2(n295), .ZN(n279) );
  INV_X1 U67 ( .A(A[11]), .ZN(n295) );
  OAI21_X1 U68 ( .B1(n276), .B2(n243), .A(n3), .ZN(n271) );
  NAND2_X1 U69 ( .A1(A[12]), .A2(n289), .ZN(n238) );
  NAND2_X1 U70 ( .A1(n287), .A2(n288), .ZN(n246) );
  INV_X1 U71 ( .A(A[12]), .ZN(n288) );
  OAI21_X1 U72 ( .B1(n269), .B2(n270), .A(n238), .ZN(n264) );
  NAND2_X1 U73 ( .A1(A[13]), .A2(n274), .ZN(n239) );
  NAND2_X1 U74 ( .A1(n272), .A2(n273), .ZN(n247) );
  INV_X1 U75 ( .A(A[13]), .ZN(n273) );
  NAND2_X1 U76 ( .A1(n257), .A2(n258), .ZN(n233) );
  INV_X1 U77 ( .A(A[15]), .ZN(n258) );
  NAND2_X1 U78 ( .A1(n265), .A2(n266), .ZN(n236) );
  INV_X1 U79 ( .A(A[14]), .ZN(n266) );
  OAI21_X1 U80 ( .B1(n263), .B2(n237), .A(n239), .ZN(n261) );
  NAND2_X1 U81 ( .A1(A[14]), .A2(n267), .ZN(n231) );
  NAND4_X1 U82 ( .A1(n233), .A2(n246), .A3(n236), .A4(n247), .ZN(n224) );
  NAND2_X1 U83 ( .A1(A[15]), .A2(n259), .ZN(n225) );
  OAI21_X1 U84 ( .B1(n249), .B2(n243), .A(n3), .ZN(n248) );
  NOR2_X1 U85 ( .A1(n250), .A2(n251), .ZN(n249) );
  NOR2_X1 U86 ( .A1(n5), .A2(n242), .ZN(n250) );
  AOI21_X1 U87 ( .B1(n230), .B2(n231), .A(n232), .ZN(n229) );
  OAI21_X1 U88 ( .B1(n234), .B2(n235), .A(n236), .ZN(n230) );
  NOR2_X1 U89 ( .A1(n243), .A2(n244), .ZN(n227) );
  NAND4_X1 U90 ( .A1(n245), .A2(n96), .A3(n98), .A4(n44), .ZN(n244) );
  NAND2_X1 U91 ( .A1(n252), .A2(n253), .ZN(n67) );
  INV_X1 U92 ( .A(A[16]), .ZN(n253) );
  NAND2_X1 U93 ( .A1(A[16]), .A2(n254), .ZN(n201) );
  NAND2_X1 U94 ( .A1(A[17]), .A2(n221), .ZN(n200) );
  NAND2_X1 U95 ( .A1(A[18]), .A2(n217), .ZN(n197) );
  NAND2_X1 U96 ( .A1(A[19]), .A2(n211), .ZN(n193) );
  NAND2_X1 U97 ( .A1(n215), .A2(n216), .ZN(n72) );
  INV_X1 U98 ( .A(A[18]), .ZN(n216) );
  NAND2_X1 U99 ( .A1(n67), .A2(n56), .ZN(n190) );
  NAND2_X1 U100 ( .A1(n219), .A2(n220), .ZN(n71) );
  INV_X1 U101 ( .A(A[17]), .ZN(n220) );
  NAND2_X1 U102 ( .A1(A[20]), .A2(n186), .ZN(n184) );
  NAND2_X1 U103 ( .A1(n165), .A2(n166), .ZN(n153) );
  INV_X1 U104 ( .A(A[23]), .ZN(n166) );
  NAND2_X1 U105 ( .A1(A[23]), .A2(n167), .ZN(n152) );
  OAI21_X1 U106 ( .B1(n175), .B2(n176), .A(n177), .ZN(n168) );
  NAND2_X1 U107 ( .A1(n173), .A2(n174), .ZN(n162) );
  INV_X1 U108 ( .A(A[22]), .ZN(n174) );
  OAI21_X1 U109 ( .B1(n112), .B2(n142), .A(n143), .ZN(n141) );
  OAI21_X1 U110 ( .B1(n134), .B2(n135), .A(n136), .ZN(n129) );
  AOI21_X1 U111 ( .B1(n120), .B2(n121), .A(n122), .ZN(n117) );
  NAND2_X1 U112 ( .A1(A[26]), .A2(n131), .ZN(n119) );
  NAND2_X1 U113 ( .A1(A[27]), .A2(n128), .ZN(n114) );
  NAND2_X1 U114 ( .A1(n139), .A2(n140), .ZN(n121) );
  INV_X1 U115 ( .A(A[25]), .ZN(n140) );
  NAND2_X1 U116 ( .A1(n146), .A2(n147), .ZN(n123) );
  INV_X1 U117 ( .A(A[24]), .ZN(n147) );
  NAND2_X1 U118 ( .A1(n126), .A2(n127), .ZN(n115) );
  INV_X1 U119 ( .A(A[27]), .ZN(n127) );
  NAND2_X1 U120 ( .A1(n132), .A2(n133), .ZN(n124) );
  INV_X1 U121 ( .A(A[26]), .ZN(n133) );
  XNOR2_X1 U122 ( .A(B[28]), .B(n352), .ZN(n109) );
  NAND2_X1 U123 ( .A1(n88), .A2(n89), .ZN(n63) );
  INV_X1 U124 ( .A(A[30]), .ZN(n89) );
  NAND2_X1 U125 ( .A1(A[29]), .A2(n100), .ZN(n92) );
  NAND2_X1 U126 ( .A1(n348), .A2(n349), .ZN(n245) );
  INV_X1 U127 ( .A(A[0]), .ZN(n349) );
  INV_X1 U128 ( .A(n353), .ZN(n351) );
  NAND2_X1 U129 ( .A1(A[0]), .A2(n350), .ZN(n204) );
  XNOR2_X1 U130 ( .A(n81), .B(n1), .ZN(SUM[31]) );
  AOI21_X1 U131 ( .B1(n63), .B2(n85), .A(n86), .ZN(n81) );
  NAND2_X1 U132 ( .A1(n101), .A2(n102), .ZN(n64) );
  INV_X1 U133 ( .A(A[29]), .ZN(n102) );
  NAND2_X1 U134 ( .A1(A[30]), .A2(n87), .ZN(n78) );
  XNOR2_X1 U135 ( .A(B[31]), .B(n352), .ZN(n82) );
  NAND2_X1 U136 ( .A1(A[31]), .A2(n84), .ZN(n75) );
  OAI21_X1 U137 ( .B1(n195), .B2(n196), .A(n197), .ZN(n194) );
  NAND4_X1 U138 ( .A1(n161), .A2(n159), .A3(n162), .A4(n153), .ZN(n55) );
  NAND2_X1 U139 ( .A1(n151), .A2(n152), .ZN(n54) );
  OAI21_X1 U140 ( .B1(n155), .B2(n156), .A(n157), .ZN(n154) );
  AOI21_X1 U141 ( .B1(n158), .B2(n159), .A(n160), .ZN(n155) );
  AND4_X1 U142 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(n7) );
  NAND2_X1 U143 ( .A1(n209), .A2(n210), .ZN(n70) );
  INV_X1 U144 ( .A(A[19]), .ZN(n210) );
  NAND2_X1 U145 ( .A1(n71), .A2(n72), .ZN(n68) );
  NAND2_X1 U146 ( .A1(A[1]), .A2(n339), .ZN(n95) );
  NAND2_X1 U147 ( .A1(n340), .A2(n341), .ZN(n96) );
  INV_X1 U148 ( .A(A[1]), .ZN(n341) );
  NAND2_X1 U149 ( .A1(n203), .A2(n204), .ZN(n97) );
  NAND2_X1 U150 ( .A1(n335), .A2(n336), .ZN(n98) );
  INV_X1 U151 ( .A(A[2]), .ZN(n336) );
  NAND2_X1 U152 ( .A1(n94), .A2(n95), .ZN(n43) );
  NAND2_X1 U153 ( .A1(n96), .A2(n97), .ZN(n94) );
  NAND2_X1 U154 ( .A1(A[2]), .A2(n334), .ZN(n42) );
  NAND2_X1 U155 ( .A1(n331), .A2(n342), .ZN(n44) );
  INV_X1 U156 ( .A(A[3]), .ZN(n342) );
  NAND2_X1 U157 ( .A1(A[3]), .A2(n330), .ZN(n45) );
  NAND2_X1 U158 ( .A1(A[4]), .A2(n320), .ZN(n34) );
  NAND2_X1 U159 ( .A1(n321), .A2(n325), .ZN(n36) );
  INV_X1 U160 ( .A(A[4]), .ZN(n325) );
  NAND2_X1 U161 ( .A1(n5), .A2(n326), .ZN(n35) );
  AND2_X1 U162 ( .A1(n98), .A2(n96), .ZN(n328) );
  NAND2_X1 U163 ( .A1(A[5]), .A2(n318), .ZN(n29) );
  NAND2_X1 U164 ( .A1(n319), .A2(n323), .ZN(n30) );
  INV_X1 U165 ( .A(A[5]), .ZN(n323) );
  NAND2_X1 U166 ( .A1(n33), .A2(n34), .ZN(n31) );
  NAND2_X1 U167 ( .A1(n35), .A2(n36), .ZN(n33) );
  NAND2_X1 U168 ( .A1(n315), .A2(n322), .ZN(n22) );
  INV_X1 U169 ( .A(A[6]), .ZN(n322) );
  OAI21_X1 U170 ( .B1(n27), .B2(n28), .A(n29), .ZN(n23) );
  NAND2_X1 U171 ( .A1(A[6]), .A2(n314), .ZN(n21) );
  NAND2_X1 U172 ( .A1(n22), .A2(n23), .ZN(n20) );
  NAND2_X1 U173 ( .A1(n310), .A2(n324), .ZN(n24) );
  INV_X1 U174 ( .A(A[7]), .ZN(n324) );
  NAND2_X1 U175 ( .A1(A[7]), .A2(n309), .ZN(n25) );
  NAND2_X1 U176 ( .A1(A[8]), .A2(n303), .ZN(n17) );
  NAND2_X1 U177 ( .A1(n304), .A2(n305), .ZN(n16) );
  INV_X1 U178 ( .A(A[8]), .ZN(n305) );
  OAI21_X1 U179 ( .B1(n306), .B2(n242), .A(n307), .ZN(n15) );
  XNOR2_X1 U180 ( .A(n10), .B(n11), .ZN(SUM[9]) );
  NAND2_X1 U181 ( .A1(n12), .A2(n13), .ZN(n10) );
  NAND2_X1 U182 ( .A1(n344), .A2(n345), .ZN(n286) );
  INV_X1 U183 ( .A(A[10]), .ZN(n345) );
  OAI21_X1 U184 ( .B1(n298), .B2(n299), .A(n13), .ZN(n293) );
  NAND2_X1 U185 ( .A1(A[10]), .A2(n346), .ZN(n283) );
  XNOR2_X1 U186 ( .A(n290), .B(n291), .ZN(SUM[11]) );
  NAND2_X1 U187 ( .A1(n278), .A2(n279), .ZN(n290) );
  OAI21_X1 U188 ( .B1(n292), .B2(n282), .A(n283), .ZN(n291) );
  XNOR2_X1 U189 ( .A(n275), .B(n271), .ZN(SUM[12]) );
  NAND2_X1 U190 ( .A1(n238), .A2(n246), .ZN(n275) );
  XNOR2_X1 U191 ( .A(n268), .B(n264), .ZN(SUM[13]) );
  NAND2_X1 U192 ( .A1(n239), .A2(n247), .ZN(n268) );
  XNOR2_X1 U193 ( .A(n262), .B(n261), .ZN(SUM[14]) );
  NAND2_X1 U194 ( .A1(n231), .A2(n236), .ZN(n262) );
  XNOR2_X1 U195 ( .A(n255), .B(n256), .ZN(SUM[15]) );
  NAND2_X1 U196 ( .A1(n225), .A2(n233), .ZN(n256) );
  NAND2_X1 U197 ( .A1(n231), .A2(n260), .ZN(n255) );
  NAND2_X1 U198 ( .A1(n261), .A2(n236), .ZN(n260) );
  OAI211_X1 U199 ( .C1(n223), .C2(n224), .A(n225), .B(n226), .ZN(n56) );
  AOI21_X1 U200 ( .B1(n227), .B2(n228), .A(n229), .ZN(n226) );
  INV_X1 U201 ( .A(n248), .ZN(n223) );
  NOR2_X1 U202 ( .A1(n240), .A2(n224), .ZN(n228) );
  NAND2_X1 U203 ( .A1(n201), .A2(n67), .ZN(n222) );
  NAND2_X1 U204 ( .A1(n190), .A2(n201), .ZN(n214) );
  NAND2_X1 U205 ( .A1(n200), .A2(n71), .ZN(n218) );
  NAND2_X1 U206 ( .A1(n213), .A2(n200), .ZN(n208) );
  NAND2_X1 U207 ( .A1(n71), .A2(n214), .ZN(n213) );
  NAND2_X1 U208 ( .A1(n197), .A2(n72), .ZN(n212) );
  OAI21_X1 U209 ( .B1(n207), .B2(n196), .A(n197), .ZN(n206) );
  NAND2_X1 U210 ( .A1(n193), .A2(n70), .ZN(n205) );
  OAI21_X1 U211 ( .B1(n190), .B2(n191), .A(n2), .ZN(n189) );
  NOR2_X1 U212 ( .A1(n183), .A2(n158), .ZN(n185) );
  OAI21_X1 U213 ( .B1(n149), .B2(n183), .A(n184), .ZN(n182) );
  NOR2_X1 U214 ( .A1(n176), .A2(n160), .ZN(n178) );
  NOR2_X1 U215 ( .A1(n156), .A2(n169), .ZN(n171) );
  XOR2_X1 U216 ( .A(n163), .B(n164), .Z(SUM[23]) );
  NAND2_X1 U217 ( .A1(n152), .A2(n153), .ZN(n164) );
  NOR2_X1 U218 ( .A1(n142), .A2(n120), .ZN(n144) );
  NOR2_X1 U219 ( .A1(n135), .A2(n122), .ZN(n137) );
  XNOR2_X1 U220 ( .A(n129), .B(n8), .ZN(SUM[26]) );
  OR2_X1 U221 ( .A1(n118), .A2(n130), .ZN(n8) );
  XNOR2_X1 U222 ( .A(n125), .B(n6), .ZN(SUM[27]) );
  AOI21_X1 U223 ( .B1(n124), .B2(n129), .A(n130), .ZN(n125) );
  OAI21_X1 U224 ( .B1(n117), .B2(n118), .A(n119), .ZN(n116) );
  NAND4_X1 U225 ( .A1(n123), .A2(n121), .A3(n124), .A4(n115), .ZN(n52) );
  OAI21_X1 U226 ( .B1(n149), .B2(n55), .A(n150), .ZN(n148) );
  NAND2_X1 U227 ( .A1(n109), .A2(n110), .ZN(n65) );
  INV_X1 U228 ( .A(A[28]), .ZN(n110) );
  NAND2_X1 U229 ( .A1(A[28]), .A2(n108), .ZN(n106) );
  OAI21_X1 U230 ( .B1(n90), .B2(n91), .A(n92), .ZN(n85) );
  OAI21_X1 U231 ( .B1(n104), .B2(n105), .A(n106), .ZN(n103) );
  XNOR2_X1 U232 ( .A(n353), .B(n347), .ZN(SUM[0]) );
  NAND2_X1 U233 ( .A1(n204), .A2(n245), .ZN(n347) );
  OAI21_X1 U234 ( .B1(n76), .B2(n77), .A(n78), .ZN(n73) );
  AOI21_X1 U235 ( .B1(n79), .B2(n64), .A(n80), .ZN(n76) );
  NAND2_X1 U236 ( .A1(n82), .A2(n83), .ZN(n62) );
  INV_X1 U237 ( .A(A[31]), .ZN(n83) );
  NAND2_X1 U238 ( .A1(n7), .A2(n50), .ZN(n49) );
  OAI21_X1 U239 ( .B1(n51), .B2(n52), .A(n4), .ZN(n50) );
  NOR2_X1 U240 ( .A1(n53), .A2(n54), .ZN(n51) );
  NOR2_X1 U241 ( .A1(n2), .A2(n55), .ZN(n53) );
  NOR2_X1 U242 ( .A1(n68), .A2(n69), .ZN(n57) );
  NOR2_X1 U243 ( .A1(n59), .A2(n60), .ZN(n58) );
  XNOR2_X1 U244 ( .A(n202), .B(n97), .ZN(SUM[1]) );
  NAND2_X1 U245 ( .A1(n96), .A2(n95), .ZN(n202) );
  XNOR2_X1 U246 ( .A(n93), .B(n43), .ZN(SUM[2]) );
  NAND2_X1 U247 ( .A1(n98), .A2(n42), .ZN(n93) );
  XNOR2_X1 U248 ( .A(n38), .B(n39), .ZN(SUM[3]) );
  NAND2_X1 U249 ( .A1(n44), .A2(n45), .ZN(n38) );
  OAI21_X1 U250 ( .B1(n40), .B2(n41), .A(n42), .ZN(n39) );
  XNOR2_X1 U251 ( .A(n37), .B(n35), .ZN(SUM[4]) );
  NAND2_X1 U252 ( .A1(n36), .A2(n34), .ZN(n37) );
  XNOR2_X1 U253 ( .A(n32), .B(n31), .ZN(SUM[5]) );
  NAND2_X1 U254 ( .A1(n30), .A2(n29), .ZN(n32) );
  XNOR2_X1 U255 ( .A(n26), .B(n23), .ZN(SUM[6]) );
  NAND2_X1 U256 ( .A1(n22), .A2(n21), .ZN(n26) );
  XNOR2_X1 U257 ( .A(n18), .B(n19), .ZN(SUM[7]) );
  NAND2_X1 U258 ( .A1(n24), .A2(n25), .ZN(n18) );
  NAND2_X1 U259 ( .A1(n20), .A2(n21), .ZN(n19) );
  XNOR2_X1 U260 ( .A(n14), .B(n15), .ZN(SUM[8]) );
  NAND2_X1 U261 ( .A1(n16), .A2(n17), .ZN(n14) );
  XNOR2_X1 U262 ( .A(n297), .B(n293), .ZN(SUM[10]) );
  NAND2_X1 U263 ( .A1(n283), .A2(n286), .ZN(n297) );
  XNOR2_X1 U264 ( .A(n218), .B(n214), .ZN(SUM[17]) );
  XNOR2_X1 U265 ( .A(n212), .B(n208), .ZN(SUM[18]) );
  XNOR2_X1 U266 ( .A(n175), .B(n178), .ZN(SUM[21]) );
  XNOR2_X1 U267 ( .A(n112), .B(n144), .ZN(SUM[24]) );
  OAI21_X1 U268 ( .B1(n112), .B2(n52), .A(n4), .ZN(n111) );
  XNOR2_X1 U269 ( .A(n85), .B(n9), .ZN(SUM[30]) );
  OR2_X1 U270 ( .A1(n77), .A2(n86), .ZN(n9) );
  NOR2_X1 U271 ( .A1(n91), .A2(n80), .ZN(n99) );
  AOI21_X1 U272 ( .B1(n62), .B2(n73), .A(n74), .ZN(n47) );
  NOR2_X1 U273 ( .A1(n105), .A2(n79), .ZN(n107) );
  INV_X1 U274 ( .A(n30), .ZN(n28) );
  INV_X1 U275 ( .A(n31), .ZN(n27) );
  INV_X1 U276 ( .A(n43), .ZN(n40) );
  XNOR2_X1 U277 ( .A(n46), .B(n351), .ZN(SUM[32]) );
  NAND3_X1 U278 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n46) );
  NAND3_X1 U279 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n48) );
  NAND2_X1 U280 ( .A1(n7), .A2(n61), .ZN(n60) );
  INV_X1 U281 ( .A(n52), .ZN(n61) );
  NAND2_X1 U282 ( .A1(n66), .A2(n67), .ZN(n59) );
  INV_X1 U283 ( .A(n55), .ZN(n66) );
  INV_X1 U284 ( .A(n70), .ZN(n69) );
  INV_X1 U285 ( .A(n75), .ZN(n74) );
  INV_X1 U286 ( .A(n82), .ZN(n84) );
  INV_X1 U287 ( .A(n78), .ZN(n86) );
  INV_X1 U288 ( .A(n88), .ZN(n87) );
  INV_X1 U289 ( .A(n63), .ZN(n77) );
  XNOR2_X1 U290 ( .A(n90), .B(n99), .ZN(SUM[29]) );
  INV_X1 U291 ( .A(n92), .ZN(n80) );
  INV_X1 U292 ( .A(n101), .ZN(n100) );
  INV_X1 U293 ( .A(n64), .ZN(n91) );
  INV_X1 U294 ( .A(n103), .ZN(n90) );
  XNOR2_X1 U295 ( .A(n104), .B(n107), .ZN(SUM[28]) );
  INV_X1 U296 ( .A(n106), .ZN(n79) );
  INV_X1 U297 ( .A(n109), .ZN(n108) );
  INV_X1 U298 ( .A(n65), .ZN(n105) );
  INV_X1 U299 ( .A(n111), .ZN(n104) );
  NAND2_X1 U300 ( .A1(n115), .A2(n116), .ZN(n113) );
  INV_X1 U301 ( .A(n126), .ZN(n128) );
  INV_X1 U302 ( .A(n119), .ZN(n130) );
  INV_X1 U303 ( .A(n132), .ZN(n131) );
  INV_X1 U304 ( .A(n124), .ZN(n118) );
  XNOR2_X1 U305 ( .A(n134), .B(n137), .ZN(SUM[25]) );
  INV_X1 U306 ( .A(n136), .ZN(n122) );
  INV_X1 U307 ( .A(n139), .ZN(n138) );
  INV_X1 U308 ( .A(n121), .ZN(n135) );
  INV_X1 U309 ( .A(n141), .ZN(n134) );
  INV_X1 U310 ( .A(n143), .ZN(n120) );
  INV_X1 U311 ( .A(n146), .ZN(n145) );
  INV_X1 U312 ( .A(n123), .ZN(n142) );
  INV_X1 U313 ( .A(n148), .ZN(n112) );
  INV_X1 U314 ( .A(n54), .ZN(n150) );
  NAND2_X1 U315 ( .A1(n153), .A2(n154), .ZN(n151) );
  INV_X1 U316 ( .A(n165), .ZN(n167) );
  AOI21_X1 U317 ( .B1(n162), .B2(n168), .A(n169), .ZN(n163) );
  XNOR2_X1 U318 ( .A(n170), .B(n171), .ZN(SUM[22]) );
  INV_X1 U319 ( .A(n157), .ZN(n169) );
  INV_X1 U320 ( .A(n173), .ZN(n172) );
  INV_X1 U321 ( .A(n162), .ZN(n156) );
  INV_X1 U322 ( .A(n168), .ZN(n170) );
  INV_X1 U323 ( .A(n177), .ZN(n160) );
  INV_X1 U324 ( .A(n180), .ZN(n179) );
  INV_X1 U325 ( .A(n159), .ZN(n176) );
  INV_X1 U326 ( .A(n182), .ZN(n175) );
  XNOR2_X1 U327 ( .A(n149), .B(n185), .ZN(SUM[20]) );
  INV_X1 U328 ( .A(n184), .ZN(n158) );
  INV_X1 U329 ( .A(n187), .ZN(n186) );
  INV_X1 U330 ( .A(n161), .ZN(n183) );
  INV_X1 U331 ( .A(n189), .ZN(n149) );
  NAND2_X1 U332 ( .A1(n70), .A2(n194), .ZN(n192) );
  INV_X1 U333 ( .A(n200), .ZN(n199) );
  INV_X1 U334 ( .A(n201), .ZN(n198) );
  NAND3_X1 U335 ( .A1(n72), .A2(n70), .A3(n71), .ZN(n191) );
  XNOR2_X1 U336 ( .A(n205), .B(n206), .ZN(SUM[19]) );
  INV_X1 U337 ( .A(n72), .ZN(n196) );
  INV_X1 U338 ( .A(n208), .ZN(n207) );
  INV_X1 U339 ( .A(n209), .ZN(n211) );
  INV_X1 U340 ( .A(n215), .ZN(n217) );
  INV_X1 U341 ( .A(n219), .ZN(n221) );
  XNOR2_X1 U342 ( .A(n222), .B(n56), .ZN(SUM[16]) );
  INV_X1 U343 ( .A(n233), .ZN(n232) );
  INV_X1 U344 ( .A(n239), .ZN(n234) );
  NAND2_X1 U345 ( .A1(n241), .A2(n352), .ZN(n240) );
  INV_X1 U346 ( .A(n242), .ZN(n241) );
  INV_X1 U347 ( .A(n252), .ZN(n254) );
  INV_X1 U348 ( .A(n257), .ZN(n259) );
  INV_X1 U349 ( .A(n247), .ZN(n237) );
  INV_X1 U350 ( .A(n264), .ZN(n263) );
  INV_X1 U351 ( .A(n265), .ZN(n267) );
  INV_X1 U352 ( .A(n246), .ZN(n270) );
  INV_X1 U353 ( .A(n271), .ZN(n269) );
  INV_X1 U354 ( .A(n272), .ZN(n274) );
  NAND2_X1 U355 ( .A1(n279), .A2(n280), .ZN(n277) );
  INV_X1 U356 ( .A(n13), .ZN(n285) );
  INV_X1 U357 ( .A(n17), .ZN(n284) );
  INV_X1 U358 ( .A(n15), .ZN(n276) );
  INV_X1 U359 ( .A(n287), .ZN(n289) );
  INV_X1 U360 ( .A(n286), .ZN(n282) );
  INV_X1 U361 ( .A(n293), .ZN(n292) );
  INV_X1 U362 ( .A(n294), .ZN(n296) );
  INV_X1 U363 ( .A(n301), .ZN(n300) );
  INV_X1 U364 ( .A(n11), .ZN(n299) );
  INV_X1 U365 ( .A(n304), .ZN(n303) );
  INV_X1 U366 ( .A(n251), .ZN(n307) );
  INV_X1 U367 ( .A(n310), .ZN(n309) );
  NAND2_X1 U368 ( .A1(n24), .A2(n311), .ZN(n308) );
  INV_X1 U369 ( .A(n315), .ZN(n314) );
  INV_X1 U370 ( .A(n22), .ZN(n313) );
  INV_X1 U371 ( .A(n29), .ZN(n317) );
  INV_X1 U372 ( .A(n319), .ZN(n318) );
  INV_X1 U373 ( .A(n34), .ZN(n316) );
  INV_X1 U374 ( .A(n321), .ZN(n320) );
  INV_X1 U375 ( .A(n35), .ZN(n306) );
  NAND3_X1 U376 ( .A1(n327), .A2(n328), .A3(n44), .ZN(n326) );
  INV_X1 U377 ( .A(n203), .ZN(n327) );
  INV_X1 U378 ( .A(n331), .ZN(n330) );
  NAND2_X1 U379 ( .A1(n44), .A2(n332), .ZN(n329) );
  INV_X1 U380 ( .A(n335), .ZN(n334) );
  INV_X1 U381 ( .A(n98), .ZN(n41) );
  INV_X1 U382 ( .A(n95), .ZN(n338) );
  INV_X1 U383 ( .A(n340), .ZN(n339) );
  INV_X1 U384 ( .A(n204), .ZN(n337) );
  INV_X1 U385 ( .A(n12), .ZN(n298) );
  INV_X1 U386 ( .A(n344), .ZN(n346) );
  INV_X1 U387 ( .A(n348), .ZN(n350) );
endmodule


module ALU_N32 ( .ALU_OPCODE({\ALU_OPCODE[6] , \ALU_OPCODE[5] , 
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), DATA1, DATA2, NEG, ZERO, CARRY, OVF, OUTALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  input \ALU_OPCODE[6] , \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] ;
  output NEG, ZERO, CARRY, OVF;
  wire   N1568, N1572, N1573, N1576, N1577, N1610, N1611, N1612, N1613, N1614,
         N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624,
         N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634,
         N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1979, N1980, N1981,
         N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991,
         N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001,
         N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011,
         \U2/U1/Z_0 , n251, n255, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n271, n272, n274, n275, n276, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n289, n291, n292, n294,
         n295, n296, n297, n298, n299, n300, n301, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n342, n343, n344, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n510, n512, n513, n514, n519, n522, n524, n526, n527, n528,
         n530, n534, n535, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n648, n649, n650,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n666, n667, n668, n669, n670, n671, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n694, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n739, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1154, n1155, n1156, n1157, n1158, n1159, n1163,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1185, n1186, n1191, n1192, n1193, n1195, n1199, n1200, n1201,
         n1204, n1205, n1206, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1239, n1240, n1241, n1242, n1243, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1339, net74079, net74084, net74087, net74089, net74092, net74095,
         net74096, net74099, net74101, net74115, net74118, net74119, net74120,
         net74121, net74123, net74124, net74128, net74130, net74133, net74135,
         net74147, net74162, net74191, net74227, net74243, net74244, net74246,
         net74249, net74263, net74287, net74292, net74295, net74296, net74299,
         net74300, net74307, net74309, net76065, net76063, net76061, net76071,
         net76069, net76067, net76091, net76089, net76087, net76107, net76149,
         net76147, net76161, net76159, net76171, net76169, net76167, net76165,
         net76163, net76177, net76479, net76488, net76487, net76493, net76501,
         net76507, net76506, net76505, net76535, net76542, net76555, net76554,
         net76553, net76566, net76573, net76578, net76759, net76778, net76781,
         net77192, net77196, net77259, net81902, net82057, net82056, net82584,
         net82652, net82651, net82724, net82738, net82899, net82925, net82924,
         net82933, net82942, net82941, net83387, net84429, net84449, net84497,
         net84496, net84507, net84505, net84530, net94830, net94964, net94951,
         net94906, net95157, n288, n287, n1207, net107648, net84501, net83745,
         n1166, n1164, n1161, net83235, n250, net83605, n249, net82884,
         net82767, n1190, n1188, n1187, n1162, n1160, net83443, net74077,
         n1170, n1169, n1168, n1167, n665, n664, n651, n647, n645, n644, n273,
         n270, n620, n362, n302, n1153, n290, net145680, net145613, net145612,
         net145611, net83422, net83343, net81160, net77211, net74076, n254,
         n252, n1172, net77228, net77226, n517, n516, n515, n511, n504,
         net84454, net83262, net82953, net82927, net82743, n501, n363, n1338,
         net94971, net94967, net84499, net83361, net82966, net82779, net112136,
         n509, n1194, n1196, n1198, n1237, n1238, n1244, n1340, n1341, n1347,
         n1348, n1349, n1351, n1352, n1353, n1354, n1357, n1358, n1359, n1361,
         n1362, n1365, n1367, n1368, n1369, n1371, n1374, n1375, n1377, n1379,
         n1383, n1388, n1390, n1391, n1392, n1393, n1395, n1398, n1399, n1401,
         n1404, n1406, n1408, n1411, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1434, n1435, n1439, n1442, n1444, n1446, n1448, n1449, n1509,
         n1511, n1517, n1520, n1527, n1528, n1530, n1535, n1536, n1537, n1538,
         n1539, n1541, n1543, n1544, n1547, n1548, n1549, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737;
  wire   [6:0] ALU_OPCODE;
  assign OUTALU[26] = net74287;
  assign OUTALU[27] = net74300;
  assign net76578 = DATA1[31];

  NOR4_X1 U259 ( .A1(n1547), .A2(n261), .A3(n262), .A4(n263), .ZN(n260) );
  NOR4_X1 U260 ( .A1(n265), .A2(n266), .A3(n267), .A4(n268), .ZN(n259) );
  NOR4_X1 U263 ( .A1(n1549), .A2(n275), .A3(n1375), .A4(n1548), .ZN(n269) );
  NOR4_X1 U265 ( .A1(n1554), .A2(n1543), .A3(n279), .A4(n280), .ZN(n278) );
  NOR4_X1 U270 ( .A1(n1559), .A2(n1539), .A3(n291), .A4(n1556), .ZN(n286) );
  OAI21_X1 U272 ( .B1(n294), .B2(n295), .A(n296), .ZN(OVF) );
  AOI22_X1 U273 ( .A1(n297), .A2(net74309), .B1(N2011), .B2(n298), .ZN(n296)
         );
  OAI21_X1 U274 ( .B1(n299), .B2(net83235), .A(n300), .ZN(n298) );
  NAND2_X1 U275 ( .A1(net84449), .A2(n301), .ZN(n300) );
  AOI21_X1 U276 ( .B1(net76573), .B2(n302), .A(n303), .ZN(n299) );
  NOR3_X1 U277 ( .A1(net74079), .A2(net83262), .A3(net76573), .ZN(n303) );
  NOR2_X1 U278 ( .A1(net76566), .A2(n304), .ZN(n297) );
  AOI22_X1 U279 ( .A1(n305), .A2(net74084), .B1(n306), .B2(n307), .ZN(n304) );
  OAI21_X1 U280 ( .B1(net76573), .B2(net74092), .A(n308), .ZN(n307) );
  AOI22_X1 U281 ( .A1(n309), .A2(n310), .B1(n252), .B2(net81160), .ZN(n308) );
  NOR2_X1 U282 ( .A1(n311), .A2(net84454), .ZN(n309) );
  AOI22_X1 U284 ( .A1(n252), .A2(net74079), .B1(n314), .B2(net84454), .ZN(n312) );
  NAND2_X1 U285 ( .A1(net76566), .A2(n315), .ZN(n295) );
  AOI22_X1 U287 ( .A1(n317), .A2(n318), .B1(n319), .B2(net74092), .ZN(n316) );
  NAND2_X1 U289 ( .A1(N2011), .A2(n320), .ZN(n318) );
  AOI22_X1 U292 ( .A1(DATA2[31]), .A2(net74263), .B1(N2010), .B2(net76578), 
        .ZN(n323) );
  OAI21_X1 U293 ( .B1(n324), .B2(net76171), .A(n325), .ZN(OUTALU[9]) );
  NAND2_X1 U294 ( .A1(n291), .A2(net76163), .ZN(n325) );
  OAI21_X1 U295 ( .B1(n281), .B2(net76171), .A(n326), .ZN(OUTALU[8]) );
  NAND2_X1 U296 ( .A1(n1554), .A2(net76165), .ZN(n326) );
  NOR4_X1 U297 ( .A1(n327), .A2(n328), .A3(n329), .A4(n330), .ZN(n324) );
  AOI21_X1 U298 ( .B1(n331), .B2(n1598), .A(n1662), .ZN(n330) );
  OAI21_X1 U299 ( .B1(n1633), .B2(n333), .A(n334), .ZN(n332) );
  AOI22_X1 U300 ( .A1(n1680), .A2(n335), .B1(n1681), .B2(n336), .ZN(n334) );
  AOI21_X1 U301 ( .B1(n337), .B2(n1682), .A(n338), .ZN(n331) );
  OAI21_X1 U302 ( .B1(n1683), .B2(n339), .A(n1555), .ZN(n338) );
  AOI21_X1 U303 ( .B1(n340), .B2(net76161), .A(n1678), .ZN(n329) );
  AOI22_X1 U304 ( .A1(DATA1[9]), .A2(net76063), .B1(net76147), .B2(n1636), 
        .ZN(n340) );
  OAI21_X1 U305 ( .B1(n1637), .B2(n1689), .A(n342), .ZN(n328) );
  AOI21_X1 U306 ( .B1(DATA1[9]), .B2(n343), .A(n344), .ZN(n342) );
  OAI21_X1 U307 ( .B1(n1417), .B2(net76493), .A(net76159), .ZN(n343) );
  NAND2_X1 U308 ( .A1(n347), .A2(n348), .ZN(n327) );
  AOI22_X1 U309 ( .A1(n349), .A2(n350), .B1(n351), .B2(n1434), .ZN(n348) );
  OR2_X1 U310 ( .A1(n353), .A2(n354), .ZN(n349) );
  OAI21_X1 U311 ( .B1(n1633), .B2(net74119), .A(n355), .ZN(n354) );
  AOI22_X1 U312 ( .A1(n1520), .A2(n335), .B1(n1517), .B2(n336), .ZN(n355) );
  OAI21_X1 U313 ( .B1(n1587), .B2(net74133), .A(n358), .ZN(n353) );
  AOI22_X1 U314 ( .A1(n359), .A2(n360), .B1(n361), .B2(n337), .ZN(n358) );
  AOI22_X1 U315 ( .A1(N1619), .A2(net76177), .B1(N1988), .B2(net76507), .ZN(
        n347) );
  OAI21_X1 U316 ( .B1(net76555), .B2(n281), .A(n364), .ZN(OUTALU[7]) );
  NAND2_X1 U317 ( .A1(net76555), .A2(n279), .ZN(n364) );
  NOR4_X1 U318 ( .A1(n365), .A2(n366), .A3(n367), .A4(n368), .ZN(n281) );
  NAND2_X1 U319 ( .A1(n369), .A2(n370), .ZN(n368) );
  AOI22_X1 U320 ( .A1(N1618), .A2(net76177), .B1(N1987), .B2(net76506), .ZN(
        n369) );
  OAI21_X1 U321 ( .B1(n1690), .B2(n371), .A(n372), .ZN(n367) );
  AOI22_X1 U322 ( .A1(n373), .A2(n374), .B1(n375), .B2(n376), .ZN(n372) );
  OAI21_X1 U323 ( .B1(n1626), .B2(n377), .A(n378), .ZN(n366) );
  AOI22_X1 U324 ( .A1(n1429), .A2(n379), .B1(n380), .B2(n381), .ZN(n378) );
  NAND2_X1 U325 ( .A1(n382), .A2(net76161), .ZN(n379) );
  AOI22_X1 U326 ( .A1(DATA1[8]), .A2(net76061), .B1(net76149), .B2(n1638), 
        .ZN(n382) );
  OAI21_X1 U327 ( .B1(n383), .B2(n1686), .A(n384), .ZN(n365) );
  AOI21_X1 U328 ( .B1(DATA1[8]), .B2(n385), .A(n386), .ZN(n384) );
  NOR3_X1 U329 ( .A1(n1683), .A2(n387), .A3(n1662), .ZN(n386) );
  OAI21_X1 U330 ( .B1(n1429), .B2(net76493), .A(net76159), .ZN(n385) );
  OAI21_X1 U331 ( .B1(n1561), .B2(net76169), .A(n389), .ZN(OUTALU[6]) );
  NAND2_X1 U332 ( .A1(n279), .A2(net76165), .ZN(n389) );
  OAI21_X1 U334 ( .B1(n394), .B2(n1653), .A(n395), .ZN(n393) );
  AOI21_X1 U335 ( .B1(n396), .B2(DATA1[7]), .A(n344), .ZN(n395) );
  OAI21_X1 U336 ( .B1(net76493), .B2(n1427), .A(net76159), .ZN(n396) );
  AOI22_X1 U337 ( .A1(n397), .A2(n398), .B1(n399), .B2(n350), .ZN(n392) );
  NAND2_X1 U338 ( .A1(n400), .A2(n401), .ZN(n399) );
  AOI21_X1 U339 ( .B1(n361), .B2(n402), .A(n403), .ZN(n401) );
  OAI21_X1 U340 ( .B1(n1575), .B2(n1687), .A(n404), .ZN(n403) );
  NAND2_X1 U341 ( .A1(n405), .A2(n406), .ZN(n404) );
  AOI22_X1 U342 ( .A1(n1520), .A2(n408), .B1(n1517), .B2(n409), .ZN(n400) );
  AOI22_X1 U343 ( .A1(n1427), .A2(n410), .B1(n411), .B2(n412), .ZN(n391) );
  OR2_X1 U344 ( .A1(n413), .A2(n414), .ZN(n412) );
  OAI21_X1 U345 ( .B1(n1605), .B2(n415), .A(n416), .ZN(n414) );
  AOI22_X1 U346 ( .A1(n1682), .A2(n402), .B1(n1680), .B2(n408), .ZN(n416) );
  OAI21_X1 U347 ( .B1(n1570), .B2(n1683), .A(n417), .ZN(n413) );
  AOI21_X1 U348 ( .B1(n1679), .B2(n406), .A(n418), .ZN(n417) );
  NAND2_X1 U349 ( .A1(n420), .A2(net76159), .ZN(n410) );
  AOI22_X1 U350 ( .A1(DATA1[7]), .A2(net76061), .B1(net76149), .B2(n1642), 
        .ZN(n420) );
  AOI22_X1 U351 ( .A1(N1617), .A2(net76177), .B1(N1986), .B2(net76505), .ZN(
        n390) );
  OAI21_X1 U352 ( .B1(n285), .B2(net76169), .A(n421), .ZN(OUTALU[5]) );
  NAND2_X1 U353 ( .A1(n280), .A2(net76163), .ZN(n421) );
  OAI21_X1 U355 ( .B1(n394), .B2(n1654), .A(n426), .ZN(n425) );
  AOI21_X1 U356 ( .B1(n427), .B2(DATA1[6]), .A(n344), .ZN(n426) );
  OAI21_X1 U357 ( .B1(net76493), .B2(n1401), .A(net76159), .ZN(n427) );
  AOI22_X1 U358 ( .A1(n397), .A2(n428), .B1(n429), .B2(n350), .ZN(n424) );
  NAND2_X1 U359 ( .A1(n430), .A2(n431), .ZN(n429) );
  AOI21_X1 U360 ( .B1(n361), .B2(n432), .A(n433), .ZN(n431) );
  OAI21_X1 U361 ( .B1(n1565), .B2(n1687), .A(n434), .ZN(n433) );
  NAND2_X1 U362 ( .A1(n405), .A2(n435), .ZN(n434) );
  AOI22_X1 U363 ( .A1(n1520), .A2(n437), .B1(n1517), .B2(n438), .ZN(n430) );
  AOI22_X1 U364 ( .A1(n1401), .A2(n439), .B1(n411), .B2(n440), .ZN(n423) );
  OR2_X1 U365 ( .A1(n441), .A2(n442), .ZN(n440) );
  OAI21_X1 U366 ( .B1(n1609), .B2(n415), .A(n443), .ZN(n442) );
  AOI22_X1 U367 ( .A1(n1682), .A2(n432), .B1(n1680), .B2(n437), .ZN(n443) );
  OAI21_X1 U368 ( .B1(n1639), .B2(n333), .A(n444), .ZN(n441) );
  AOI21_X1 U369 ( .B1(n445), .B2(n446), .A(n418), .ZN(n444) );
  NAND2_X1 U370 ( .A1(n447), .A2(net76159), .ZN(n439) );
  AOI22_X1 U371 ( .A1(DATA1[6]), .A2(net76061), .B1(net76149), .B2(n1643), 
        .ZN(n447) );
  AOI22_X1 U372 ( .A1(N1616), .A2(net76177), .B1(N1985), .B2(net76507), .ZN(
        n422) );
  OAI21_X1 U373 ( .B1(net76554), .B2(n285), .A(n448), .ZN(OUTALU[4]) );
  NAND2_X1 U374 ( .A1(net76554), .A2(n282), .ZN(n448) );
  NOR3_X1 U375 ( .A1(n449), .A2(n450), .A3(n451), .ZN(n285) );
  OAI21_X1 U376 ( .B1(n1648), .B2(n1689), .A(n452), .ZN(n451) );
  OAI21_X1 U377 ( .B1(n453), .B2(n454), .A(n350), .ZN(n452) );
  OAI21_X1 U378 ( .B1(n1633), .B2(n1692), .A(n455), .ZN(n454) );
  AOI22_X1 U379 ( .A1(n1517), .A2(n335), .B1(n456), .B2(n336), .ZN(n455) );
  NAND2_X1 U380 ( .A1(n457), .A2(n458), .ZN(n453) );
  AOI22_X1 U381 ( .A1(n459), .A2(n1442), .B1(n359), .B2(n460), .ZN(n458) );
  NOR2_X1 U382 ( .A1(n1576), .A2(n1693), .ZN(n459) );
  AOI22_X1 U383 ( .A1(n1520), .A2(n337), .B1(n405), .B2(n461), .ZN(n457) );
  OAI21_X1 U384 ( .B1(n462), .B2(n394), .A(n463), .ZN(n450) );
  AOI21_X1 U385 ( .B1(DATA1[5]), .B2(n464), .A(n344), .ZN(n463) );
  OAI21_X1 U386 ( .B1(n1425), .B2(net76493), .A(net76159), .ZN(n464) );
  NAND2_X1 U387 ( .A1(n465), .A2(n1434), .ZN(n394) );
  NAND2_X1 U388 ( .A1(n466), .A2(n467), .ZN(n449) );
  AOI22_X1 U389 ( .A1(n1425), .A2(n468), .B1(n411), .B2(n469), .ZN(n467) );
  NAND2_X1 U390 ( .A1(n470), .A2(n471), .ZN(n469) );
  AOI21_X1 U391 ( .B1(n461), .B2(n1679), .A(n1612), .ZN(n471) );
  AOI22_X1 U392 ( .A1(n1680), .A2(n337), .B1(n1681), .B2(n335), .ZN(n472) );
  AOI21_X1 U393 ( .B1(n473), .B2(n1682), .A(n474), .ZN(n470) );
  OAI21_X1 U394 ( .B1(n1683), .B2(n475), .A(n1555), .ZN(n474) );
  NAND2_X1 U395 ( .A1(n476), .A2(net76159), .ZN(n468) );
  AOI22_X1 U396 ( .A1(DATA1[5]), .A2(net76061), .B1(net76149), .B2(n1646), 
        .ZN(n476) );
  AOI22_X1 U397 ( .A1(N1615), .A2(net76177), .B1(N1984), .B2(net76506), .ZN(
        n466) );
  OAI21_X1 U398 ( .B1(n1552), .B2(net76169), .A(n477), .ZN(OUTALU[3]) );
  NAND2_X1 U399 ( .A1(n282), .A2(net76163), .ZN(n477) );
  NOR3_X1 U401 ( .A1(n482), .A2(n483), .A3(n484), .ZN(n481) );
  OAI33_X1 U402 ( .A1(n485), .A2(n1439), .A3(n1690), .B1(n1683), .B2(n486), 
        .B3(n1662), .ZN(n484) );
  NOR2_X1 U403 ( .A1(n487), .A2(n1651), .ZN(n483) );
  AOI21_X1 U404 ( .B1(net76149), .B2(n1687), .A(net76488), .ZN(n487) );
  OAI21_X1 U405 ( .B1(n1635), .B2(n377), .A(n489), .ZN(n482) );
  AOI22_X1 U406 ( .A1(n1442), .A2(n490), .B1(n380), .B2(n491), .ZN(n489) );
  OAI21_X1 U407 ( .B1(n1662), .B2(n492), .A(n493), .ZN(n380) );
  NAND2_X1 U408 ( .A1(n1520), .A2(n350), .ZN(n493) );
  NAND2_X1 U409 ( .A1(n494), .A2(n495), .ZN(n490) );
  AOI22_X1 U410 ( .A1(n1541), .A2(n350), .B1(n1449), .B2(net76065), .ZN(n495)
         );
  AOI21_X1 U411 ( .B1(net76149), .B2(n1651), .A(net76488), .ZN(n494) );
  AOI21_X1 U412 ( .B1(n411), .B2(n1682), .A(n497), .ZN(n377) );
  NOR2_X1 U413 ( .A1(n1692), .A2(n1701), .ZN(n497) );
  AOI21_X1 U414 ( .B1(N1983), .B2(net76506), .A(n1560), .ZN(n480) );
  AOI21_X1 U415 ( .B1(n418), .B2(n411), .A(n344), .ZN(n370) );
  NAND2_X1 U416 ( .A1(N1614), .A2(net76177), .ZN(n479) );
  AOI22_X1 U417 ( .A1(n373), .A2(n381), .B1(n375), .B2(n498), .ZN(n478) );
  OAI21_X1 U418 ( .B1(n333), .B2(n1662), .A(net74120), .ZN(n375) );
  OAI21_X1 U419 ( .B1(n1662), .B2(n415), .A(n499), .ZN(n373) );
  NAND2_X1 U420 ( .A1(n1517), .A2(n350), .ZN(n499) );
  OAI21_X1 U443 ( .B1(n1551), .B2(net76169), .A(n538), .ZN(OUTALU[2]) );
  NAND2_X1 U444 ( .A1(n283), .A2(net76165), .ZN(n538) );
  NOR3_X1 U446 ( .A1(n543), .A2(n544), .A3(n545), .ZN(n542) );
  NOR3_X1 U447 ( .A1(n546), .A2(n547), .A3(n1687), .ZN(n545) );
  NOR2_X1 U448 ( .A1(n548), .A2(n1652), .ZN(n543) );
  AOI21_X1 U449 ( .B1(net76149), .B2(n1694), .A(net76488), .ZN(n548) );
  AOI21_X1 U450 ( .B1(n388), .B2(n1354), .A(n549), .ZN(n541) );
  AOI21_X1 U451 ( .B1(n550), .B2(n551), .A(n552), .ZN(n549) );
  AOI21_X1 U452 ( .B1(n1509), .B2(n406), .A(n553), .ZN(n551) );
  NOR2_X1 U453 ( .A1(n554), .A2(net74115), .ZN(n553) );
  NOR4_X1 U454 ( .A1(n555), .A2(n556), .A3(n557), .A4(n558), .ZN(n554) );
  NOR2_X1 U455 ( .A1(n1704), .A2(n1646), .ZN(n558) );
  NAND2_X1 U456 ( .A1(n559), .A2(n560), .ZN(n406) );
  AOI22_X1 U457 ( .A1(DATA1[7]), .A2(net76067), .B1(DATA1[6]), .B2(n1530), 
        .ZN(n560) );
  AOI22_X1 U458 ( .A1(DATA1[9]), .A2(net76087), .B1(DATA1[8]), .B2(net76781), 
        .ZN(n559) );
  AOI22_X1 U459 ( .A1(n562), .A2(n402), .B1(n563), .B2(n408), .ZN(n550) );
  AOI22_X1 U460 ( .A1(n1439), .A2(n565), .B1(net76501), .B2(n566), .ZN(n540)
         );
  NAND2_X1 U461 ( .A1(n567), .A2(net76159), .ZN(n565) );
  AOI22_X1 U462 ( .A1(n1448), .A2(net76061), .B1(net76149), .B2(n1652), .ZN(
        n567) );
  AOI22_X1 U463 ( .A1(N1613), .A2(net76177), .B1(N1982), .B2(net76505), .ZN(
        n539) );
  OAI21_X1 U464 ( .B1(net74296), .B2(net76167), .A(n568), .ZN(OUTALU[29]) );
  NAND2_X1 U465 ( .A1(n284), .A2(net76165), .ZN(n568) );
  AOI21_X1 U467 ( .B1(DATA1[30]), .B2(n573), .A(n574), .ZN(n572) );
  OAI21_X1 U468 ( .B1(n1664), .B2(n575), .A(n1544), .ZN(n574) );
  NAND2_X1 U469 ( .A1(n576), .A2(n577), .ZN(n575) );
  OAI21_X1 U470 ( .B1(DATA2[30]), .B2(net76493), .A(net76159), .ZN(n573) );
  AOI22_X1 U471 ( .A1(n534), .A2(n578), .B1(DATA2[30]), .B2(n579), .ZN(n571)
         );
  NAND2_X1 U472 ( .A1(n580), .A2(net76159), .ZN(n579) );
  AOI22_X1 U473 ( .A1(DATA1[30]), .A2(net76061), .B1(net76149), .B2(net74249), 
        .ZN(n580) );
  AOI22_X1 U474 ( .A1(n581), .A2(n582), .B1(n1430), .B2(net74095), .ZN(n570)
         );
  NAND2_X1 U475 ( .A1(n583), .A2(n584), .ZN(n581) );
  NOR3_X1 U476 ( .A1(n585), .A2(n586), .A3(n587), .ZN(n584) );
  AOI21_X1 U478 ( .B1(n589), .B2(n590), .A(net74119), .ZN(n586) );
  AOI22_X1 U480 ( .A1(DATA1[27]), .A2(net76089), .B1(net76781), .B2(DATA1[28]), 
        .ZN(n589) );
  AOI22_X1 U482 ( .A1(n1517), .A2(n593), .B1(n1442), .B2(n594), .ZN(n583) );
  AOI22_X1 U483 ( .A1(N1640), .A2(net76177), .B1(N2009), .B2(net76507), .ZN(
        n569) );
  OAI21_X1 U484 ( .B1(n1374), .B2(net76167), .A(n595), .ZN(OUTALU[28]) );
  NAND2_X1 U485 ( .A1(n271), .A2(net76165), .ZN(n595) );
  AOI21_X1 U487 ( .B1(n600), .B2(n360), .A(n601), .ZN(n599) );
  OAI21_X1 U488 ( .B1(net74115), .B2(n1664), .A(net74120), .ZN(n600) );
  NOR2_X1 U489 ( .A1(net74119), .A2(n1701), .ZN(n534) );
  AOI22_X1 U490 ( .A1(DATA1[29]), .A2(n602), .B1(DATA2[29]), .B2(n603), .ZN(
        n598) );
  NAND2_X1 U491 ( .A1(n604), .A2(net76161), .ZN(n603) );
  AOI22_X1 U492 ( .A1(DATA1[29]), .A2(net76061), .B1(net76149), .B2(net74246), 
        .ZN(n604) );
  OAI21_X1 U493 ( .B1(DATA2[29]), .B2(net76493), .A(net76159), .ZN(n602) );
  AOI22_X1 U494 ( .A1(n605), .A2(n582), .B1(n1428), .B2(net74095), .ZN(n597)
         );
  OR2_X1 U495 ( .A1(n606), .A2(n607), .ZN(n605) );
  OAI21_X1 U496 ( .B1(n1628), .B2(net74133), .A(n608), .ZN(n607) );
  AOI22_X1 U497 ( .A1(n1520), .A2(n609), .B1(n1517), .B2(n610), .ZN(n608) );
  NAND2_X1 U498 ( .A1(n612), .A2(n613), .ZN(n606) );
  AOI21_X1 U499 ( .B1(n1442), .B2(n614), .A(n615), .ZN(n613) );
  AOI21_X1 U500 ( .B1(n616), .B2(n617), .A(net74119), .ZN(n615) );
  AOI22_X1 U501 ( .A1(DATA1[28]), .A2(net76067), .B1(n1527), .B2(DATA1[29]), 
        .ZN(n617) );
  AOI22_X1 U502 ( .A1(DATA1[26]), .A2(net76089), .B1(DATA1[27]), .B2(net76781), 
        .ZN(n616) );
  AOI22_X1 U503 ( .A1(n359), .A2(n346), .B1(n361), .B2(n618), .ZN(n612) );
  AOI22_X1 U504 ( .A1(N1639), .A2(net76177), .B1(N2008), .B2(net76506), .ZN(
        n596) );
  AOI21_X1 U507 ( .B1(DATA1[28]), .B2(n624), .A(n625), .ZN(n623) );
  OAI21_X1 U508 ( .B1(net74115), .B2(n626), .A(n1544), .ZN(n625) );
  NOR2_X1 U509 ( .A1(net74295), .A2(net74101), .ZN(n601) );
  OR2_X1 U510 ( .A1(n1583), .A2(n627), .ZN(n626) );
  OAI21_X1 U511 ( .B1(DATA2[28]), .B2(net76493), .A(net76159), .ZN(n624) );
  AOI22_X1 U512 ( .A1(n628), .A2(n519), .B1(DATA2[28]), .B2(n629), .ZN(n622)
         );
  NAND2_X1 U513 ( .A1(n630), .A2(net76159), .ZN(n629) );
  AOI22_X1 U514 ( .A1(DATA1[28]), .A2(net76061), .B1(net76149), .B2(net74243), 
        .ZN(n630) );
  AOI22_X1 U515 ( .A1(n631), .A2(n582), .B1(n1424), .B2(net74095), .ZN(n621)
         );
  OR2_X1 U516 ( .A1(n632), .A2(n633), .ZN(n631) );
  OAI21_X1 U517 ( .B1(n1594), .B2(n1692), .A(n634), .ZN(n633) );
  AOI22_X1 U518 ( .A1(n1517), .A2(n635), .B1(n456), .B2(n636), .ZN(n634) );
  NAND2_X1 U519 ( .A1(n637), .A2(n638), .ZN(n632) );
  AOI21_X1 U520 ( .B1(n359), .B2(n639), .A(n640), .ZN(n638) );
  NOR3_X1 U521 ( .A1(n485), .A2(n1694), .A3(n1687), .ZN(n640) );
  AOI22_X1 U522 ( .A1(n405), .A2(n641), .B1(n1520), .B2(n642), .ZN(n637) );
  OAI21_X1 U528 ( .B1(n652), .B2(n1688), .A(n653), .ZN(n649) );
  OAI21_X1 U529 ( .B1(n654), .B2(net76488), .A(DATA1[27]), .ZN(n653) );
  NOR2_X1 U530 ( .A1(DATA2[27]), .A2(net76493), .ZN(n654) );
  NAND2_X1 U531 ( .A1(n655), .A2(n656), .ZN(n648) );
  AOI22_X1 U532 ( .A1(net74130), .A2(n657), .B1(n658), .B2(n659), .ZN(n656) );
  AOI22_X1 U533 ( .A1(DATA2[27]), .A2(n660), .B1(n661), .B2(n662), .ZN(n655)
         );
  NAND2_X1 U534 ( .A1(n663), .A2(net76159), .ZN(n660) );
  AOI22_X1 U535 ( .A1(DATA1[27]), .A2(net76061), .B1(net76149), .B2(n1586), 
        .ZN(n663) );
  NAND2_X1 U541 ( .A1(n667), .A2(n668), .ZN(n513) );
  AOI22_X1 U542 ( .A1(DATA1[26]), .A2(net76067), .B1(DATA1[27]), .B2(n1527), 
        .ZN(n668) );
  AOI22_X1 U543 ( .A1(DATA1[24]), .A2(net76087), .B1(DATA1[25]), .B2(net76781), 
        .ZN(n667) );
  OAI21_X1 U544 ( .B1(n276), .B2(net76167), .A(n669), .ZN(OUTALU[25]) );
  NAND2_X1 U545 ( .A1(n274), .A2(net76165), .ZN(n669) );
  NOR4_X1 U547 ( .A1(n674), .A2(n675), .A3(n650), .A4(n676), .ZN(n673) );
  NOR3_X1 U548 ( .A1(net74128), .A2(n1585), .A3(net74115), .ZN(n676) );
  OAI21_X1 U549 ( .B1(n1566), .B2(n1688), .A(n677), .ZN(n675) );
  OAI21_X1 U550 ( .B1(n678), .B2(net76488), .A(DATA1[26]), .ZN(n677) );
  NOR2_X1 U551 ( .A1(DATA2[26]), .A2(net76493), .ZN(n678) );
  NOR2_X1 U552 ( .A1(net74128), .A2(n1695), .ZN(n628) );
  NAND2_X1 U553 ( .A1(n679), .A2(n680), .ZN(n674) );
  AOI22_X1 U554 ( .A1(net74130), .A2(n681), .B1(n658), .B2(n682), .ZN(n680) );
  AOI22_X1 U555 ( .A1(DATA2[26]), .A2(n683), .B1(n661), .B2(n1562), .ZN(n679)
         );
  NAND2_X1 U556 ( .A1(n685), .A2(net76159), .ZN(n683) );
  AOI22_X1 U557 ( .A1(DATA1[26]), .A2(net76063), .B1(net76149), .B2(n1588), 
        .ZN(n685) );
  OAI21_X1 U559 ( .B1(n510), .B2(n1677), .A(n687), .ZN(n686) );
  NAND2_X1 U560 ( .A1(N1636), .A2(net76177), .ZN(n687) );
  AOI22_X1 U561 ( .A1(net74123), .A2(n688), .B1(net74124), .B2(n593), .ZN(n671) );
  AOI22_X1 U562 ( .A1(n512), .A2(n592), .B1(net76501), .B2(n588), .ZN(n670) );
  NAND2_X1 U563 ( .A1(n689), .A2(n690), .ZN(n588) );
  AOI21_X1 U564 ( .B1(DATA1[25]), .B2(net76069), .A(n691), .ZN(n690) );
  AOI22_X1 U565 ( .A1(DATA1[26]), .A2(n1527), .B1(DATA1[24]), .B2(net76781), 
        .ZN(n689) );
  OAI21_X1 U566 ( .B1(net76553), .B2(n276), .A(n692), .ZN(OUTALU[24]) );
  NAND2_X1 U567 ( .A1(net76555), .A2(n275), .ZN(n692) );
  OAI21_X1 U569 ( .B1(net74162), .B2(n1590), .A(n697), .ZN(n696) );
  AOI22_X1 U570 ( .A1(n1417), .A2(net74095), .B1(N1635), .B2(net76177), .ZN(
        n697) );
  AOI22_X1 U572 ( .A1(net74123), .A2(n611), .B1(net74124), .B2(n610), .ZN(n699) );
  AOI22_X1 U573 ( .A1(net76479), .A2(n609), .B1(n514), .B2(n618), .ZN(n698) );
  NAND2_X1 U574 ( .A1(n700), .A2(n701), .ZN(n618) );
  AOI22_X1 U575 ( .A1(DATA1[24]), .A2(net76067), .B1(DATA1[25]), .B2(n1528), 
        .ZN(n701) );
  AOI22_X1 U576 ( .A1(DATA1[22]), .A2(net76087), .B1(DATA1[23]), .B2(net76781), 
        .ZN(n700) );
  OAI21_X1 U577 ( .B1(n339), .B2(n1664), .A(n702), .ZN(n694) );
  AOI22_X1 U578 ( .A1(n703), .A2(n704), .B1(DATA2[25]), .B2(n705), .ZN(n702)
         );
  NAND2_X1 U579 ( .A1(n706), .A2(net76161), .ZN(n705) );
  AOI22_X1 U580 ( .A1(DATA1[25]), .A2(net76063), .B1(net76147), .B2(n1591), 
        .ZN(n706) );
  NOR2_X1 U581 ( .A1(n704), .A2(n707), .ZN(n339) );
  OAI21_X1 U582 ( .B1(n1576), .B2(n1695), .A(n708), .ZN(n704) );
  NAND2_X1 U583 ( .A1(net76542), .A2(n460), .ZN(n708) );
  AOI21_X1 U585 ( .B1(DATA1[25]), .B2(n711), .A(n650), .ZN(n710) );
  OAI21_X1 U586 ( .B1(DATA2[25]), .B2(net76493), .A(net76159), .ZN(n711) );
  AOI22_X1 U587 ( .A1(net74130), .A2(n351), .B1(n658), .B2(n346), .ZN(n709) );
  OAI21_X1 U588 ( .B1(n1648), .B2(n1695), .A(n712), .ZN(n351) );
  NAND2_X1 U589 ( .A1(n562), .A2(n1656), .ZN(n712) );
  OAI21_X1 U590 ( .B1(n714), .B2(net76167), .A(n715), .ZN(OUTALU[23]) );
  NAND2_X1 U591 ( .A1(n275), .A2(net76165), .ZN(n715) );
  NAND2_X1 U592 ( .A1(n716), .A2(n717), .ZN(n275) );
  NOR4_X1 U593 ( .A1(n718), .A2(n719), .A3(n720), .A4(n721), .ZN(n717) );
  AOI21_X1 U594 ( .B1(n722), .B2(net76161), .A(n1668), .ZN(n721) );
  AOI22_X1 U595 ( .A1(DATA1[24]), .A2(net76063), .B1(net76147), .B2(n1593), 
        .ZN(n722) );
  NOR2_X1 U596 ( .A1(n371), .A2(n713), .ZN(n720) );
  AOI21_X1 U597 ( .B1(n562), .B2(n723), .A(n1641), .ZN(n371) );
  AOI22_X1 U598 ( .A1(net76542), .A2(n639), .B1(n465), .B2(n725), .ZN(n724) );
  OAI21_X1 U599 ( .B1(n726), .B2(n1593), .A(net74292), .ZN(n719) );
  AOI21_X1 U600 ( .B1(net76149), .B2(n1668), .A(net76488), .ZN(n726) );
  OAI21_X1 U601 ( .B1(n1623), .B2(n522), .A(n727), .ZN(n718) );
  AOI22_X1 U602 ( .A1(n661), .A2(n1564), .B1(net74123), .B2(n636), .ZN(n727)
         );
  NOR2_X1 U603 ( .A1(n728), .A2(n707), .ZN(n387) );
  NOR2_X1 U604 ( .A1(n729), .A2(n730), .ZN(n716) );
  AOI22_X1 U606 ( .A1(n1429), .A2(net74095), .B1(N1634), .B2(net76177), .ZN(
        n731) );
  OAI21_X1 U607 ( .B1(n383), .B2(net74128), .A(n732), .ZN(n729) );
  AOI22_X1 U608 ( .A1(net76479), .A2(n642), .B1(net76501), .B2(n733), .ZN(n732) );
  AOI21_X1 U609 ( .B1(n562), .B2(n519), .A(n728), .ZN(n383) );
  OAI21_X1 U610 ( .B1(n1583), .B2(n1695), .A(n734), .ZN(n728) );
  NAND2_X1 U611 ( .A1(net76542), .A2(n735), .ZN(n734) );
  OAI21_X1 U612 ( .B1(n736), .B2(net76167), .A(n737), .ZN(OUTALU[22]) );
  NAND2_X1 U613 ( .A1(n1375), .A2(net76165), .ZN(n737) );
  OAI21_X1 U615 ( .B1(net74162), .B2(n1595), .A(n742), .ZN(n741) );
  AOI22_X1 U616 ( .A1(n1427), .A2(net74095), .B1(N1633), .B2(net76177), .ZN(
        n742) );
  AOI22_X1 U618 ( .A1(net74124), .A2(n666), .B1(n512), .B2(n524), .ZN(n744) );
  AOI22_X1 U619 ( .A1(net76501), .A2(n530), .B1(n703), .B2(n407), .ZN(n743) );
  OAI21_X1 U620 ( .B1(n652), .B2(n1693), .A(n1584), .ZN(n407) );
  NAND2_X1 U621 ( .A1(n745), .A2(n746), .ZN(n530) );
  AOI22_X1 U622 ( .A1(DATA1[22]), .A2(net76067), .B1(DATA1[23]), .B2(n1527), 
        .ZN(n746) );
  AOI22_X1 U623 ( .A1(DATA1[20]), .A2(net76087), .B1(DATA1[21]), .B2(net76781), 
        .ZN(n745) );
  OAI21_X1 U624 ( .B1(n1632), .B2(n747), .A(n748), .ZN(n739) );
  AOI22_X1 U625 ( .A1(DATA2[23]), .A2(n749), .B1(n661), .B2(n419), .ZN(n748)
         );
  NAND2_X1 U626 ( .A1(n750), .A2(n1584), .ZN(n419) );
  OAI21_X1 U627 ( .B1(net74244), .B2(n1695), .A(n752), .ZN(n751) );
  NAND2_X1 U628 ( .A1(net76542), .A2(n753), .ZN(n752) );
  AOI21_X1 U629 ( .B1(n562), .B2(n1578), .A(n754), .ZN(n750) );
  NAND2_X1 U630 ( .A1(n755), .A2(net76159), .ZN(n749) );
  AOI22_X1 U631 ( .A1(DATA1[23]), .A2(net76063), .B1(net76147), .B2(n1599), 
        .ZN(n755) );
  AOI21_X1 U633 ( .B1(DATA1[23]), .B2(n758), .A(n650), .ZN(n757) );
  OAI21_X1 U634 ( .B1(DATA2[23]), .B2(net76493), .A(net76159), .ZN(n758) );
  AOI22_X1 U635 ( .A1(n759), .A2(n566), .B1(n658), .B2(n398), .ZN(n756) );
  OAI21_X1 U636 ( .B1(n264), .B2(net76169), .A(n760), .ZN(OUTALU[21]) );
  NAND2_X1 U637 ( .A1(n1548), .A2(net76167), .ZN(n760) );
  NOR4_X1 U638 ( .A1(n761), .A2(n762), .A3(n763), .A4(n764), .ZN(n736) );
  OAI21_X1 U639 ( .B1(net74162), .B2(n1600), .A(n765), .ZN(n764) );
  AOI22_X1 U640 ( .A1(n1401), .A2(net74095), .B1(N1632), .B2(net76177), .ZN(
        n765) );
  NAND2_X1 U641 ( .A1(n766), .A2(n767), .ZN(n763) );
  AOI22_X1 U642 ( .A1(net74124), .A2(n688), .B1(n512), .B2(n593), .ZN(n767) );
  AOI22_X1 U643 ( .A1(n514), .A2(n592), .B1(n703), .B2(n436), .ZN(n766) );
  OAI21_X1 U644 ( .B1(n1566), .B2(n1693), .A(n768), .ZN(n436) );
  NAND2_X1 U645 ( .A1(n769), .A2(n770), .ZN(n592) );
  AOI22_X1 U646 ( .A1(DATA1[21]), .A2(net76067), .B1(DATA1[22]), .B2(n1528), 
        .ZN(n770) );
  AOI22_X1 U647 ( .A1(DATA1[19]), .A2(net76087), .B1(DATA1[20]), .B2(net76781), 
        .ZN(n769) );
  OAI21_X1 U648 ( .B1(n1634), .B2(n747), .A(n771), .ZN(n762) );
  AOI22_X1 U649 ( .A1(DATA2[22]), .A2(n772), .B1(n661), .B2(n446), .ZN(n771)
         );
  NAND2_X1 U650 ( .A1(n773), .A2(n768), .ZN(n446) );
  AOI21_X1 U651 ( .B1(n774), .B2(n1509), .A(n775), .ZN(n768) );
  AOI21_X1 U653 ( .B1(n562), .B2(n577), .A(n754), .ZN(n773) );
  NAND2_X1 U654 ( .A1(n777), .A2(net76161), .ZN(n772) );
  AOI22_X1 U655 ( .A1(DATA1[22]), .A2(net76063), .B1(net76149), .B2(n1601), 
        .ZN(n777) );
  NAND2_X1 U656 ( .A1(n778), .A2(n779), .ZN(n761) );
  AOI21_X1 U657 ( .B1(DATA1[22]), .B2(n780), .A(n650), .ZN(n779) );
  OAI21_X1 U658 ( .B1(DATA2[22]), .B2(net76493), .A(net76161), .ZN(n780) );
  AOI22_X1 U659 ( .A1(n759), .A2(n781), .B1(n658), .B2(n428), .ZN(n778) );
  OAI21_X1 U660 ( .B1(net76553), .B2(n264), .A(n782), .ZN(OUTALU[20]) );
  NAND2_X1 U661 ( .A1(net76554), .A2(n262), .ZN(n782) );
  NOR4_X1 U662 ( .A1(n783), .A2(n784), .A3(n785), .A4(n786), .ZN(n264) );
  OAI21_X1 U663 ( .B1(net74162), .B2(n1603), .A(n787), .ZN(n786) );
  AOI22_X1 U664 ( .A1(n1425), .A2(net74095), .B1(N1631), .B2(net76177), .ZN(
        n787) );
  NAND2_X1 U665 ( .A1(n788), .A2(n789), .ZN(n785) );
  AOI22_X1 U666 ( .A1(net74123), .A2(n346), .B1(net74124), .B2(n611), .ZN(n789) );
  AOI22_X1 U667 ( .A1(net76479), .A2(n610), .B1(net76501), .B2(n609), .ZN(n788) );
  NAND2_X1 U668 ( .A1(n790), .A2(n791), .ZN(n609) );
  AOI22_X1 U669 ( .A1(DATA1[20]), .A2(net76067), .B1(DATA1[21]), .B2(n1527), 
        .ZN(n791) );
  AOI22_X1 U670 ( .A1(DATA1[18]), .A2(net76089), .B1(DATA1[19]), .B2(net76781), 
        .ZN(n790) );
  OAI21_X1 U671 ( .B1(n475), .B2(n1664), .A(n792), .ZN(n784) );
  AOI22_X1 U672 ( .A1(n703), .A2(n793), .B1(DATA2[21]), .B2(n794), .ZN(n792)
         );
  NAND2_X1 U673 ( .A1(n795), .A2(net76159), .ZN(n794) );
  AOI22_X1 U674 ( .A1(DATA1[21]), .A2(net76063), .B1(net76149), .B2(n1604), 
        .ZN(n795) );
  NOR2_X1 U675 ( .A1(n793), .A2(n754), .ZN(n475) );
  OAI21_X1 U676 ( .B1(n1597), .B2(net74115), .A(n796), .ZN(n793) );
  AOI22_X1 U677 ( .A1(n562), .A2(n360), .B1(n1509), .B2(n460), .ZN(n796) );
  NAND2_X1 U678 ( .A1(n797), .A2(n798), .ZN(n783) );
  AOI21_X1 U679 ( .B1(DATA1[21]), .B2(n799), .A(n650), .ZN(n798) );
  OAI21_X1 U680 ( .B1(DATA2[21]), .B2(net76493), .A(net76161), .ZN(n799) );
  AOI22_X1 U681 ( .A1(n759), .A2(n1656), .B1(n658), .B2(n800), .ZN(n797) );
  NOR2_X1 U682 ( .A1(net74135), .A2(n1700), .ZN(n759) );
  AOI22_X1 U683 ( .A1(n261), .A2(net76163), .B1(net76554), .B2(n268), .ZN(n801) );
  NOR3_X1 U685 ( .A1(n806), .A2(n544), .A3(n807), .ZN(n805) );
  NOR3_X1 U686 ( .A1(n546), .A2(n808), .A3(n1687), .ZN(n807) );
  NOR2_X1 U687 ( .A1(n809), .A2(n1655), .ZN(n806) );
  AOI21_X1 U688 ( .B1(net76149), .B2(n1696), .A(net76488), .ZN(n809) );
  AOI21_X1 U689 ( .B1(n388), .B2(n1567), .A(n810), .ZN(n804) );
  AOI21_X1 U690 ( .B1(n811), .B2(n812), .A(n552), .ZN(n810) );
  AOI21_X1 U691 ( .B1(n1687), .B2(n1665), .A(n703), .ZN(n552) );
  AOI22_X1 U692 ( .A1(n576), .A2(n813), .B1(n465), .B2(n435), .ZN(n812) );
  NAND2_X1 U693 ( .A1(n814), .A2(n815), .ZN(n435) );
  AOI22_X1 U694 ( .A1(DATA1[6]), .A2(net76067), .B1(DATA1[5]), .B2(n1527), 
        .ZN(n815) );
  AOI22_X1 U695 ( .A1(DATA1[8]), .A2(net76089), .B1(DATA1[7]), .B2(net76781), 
        .ZN(n814) );
  NAND2_X1 U696 ( .A1(n816), .A2(n817), .ZN(n813) );
  AOI21_X1 U697 ( .B1(n1446), .B2(net76071), .A(n818), .ZN(n817) );
  AOI22_X1 U698 ( .A1(n1449), .A2(net76089), .B1(n1448), .B2(net76781), .ZN(
        n816) );
  AOI22_X1 U699 ( .A1(n1511), .A2(n432), .B1(n563), .B2(n437), .ZN(n811) );
  NOR2_X1 U700 ( .A1(n1687), .A2(n1701), .ZN(n388) );
  AOI22_X1 U701 ( .A1(DATA2[2]), .A2(n820), .B1(net76501), .B2(n781), .ZN(n803) );
  NAND2_X1 U702 ( .A1(n821), .A2(net76159), .ZN(n820) );
  AOI22_X1 U703 ( .A1(n1446), .A2(net76063), .B1(net76147), .B2(n1655), .ZN(
        n821) );
  AOI22_X1 U704 ( .A1(N1612), .A2(net76177), .B1(N1981), .B2(net76507), .ZN(
        n802) );
  AOI22_X1 U705 ( .A1(n262), .A2(net76163), .B1(net76555), .B2(n263), .ZN(n822) );
  NAND2_X1 U706 ( .A1(n823), .A2(n824), .ZN(n262) );
  NOR4_X1 U707 ( .A1(n825), .A2(n1607), .A3(n650), .A4(n826), .ZN(n824) );
  NOR3_X1 U708 ( .A1(n713), .A2(n1439), .A3(n485), .ZN(n826) );
  NAND2_X1 U709 ( .A1(n1442), .A2(n582), .ZN(n713) );
  AOI21_X1 U710 ( .B1(n828), .B2(DATA1[20]), .A(n1608), .ZN(n827) );
  OAI21_X1 U711 ( .B1(net76487), .B2(n830), .A(DATA2[20]), .ZN(n829) );
  OAI21_X1 U712 ( .B1(DATA1[20]), .B2(net76493), .A(n831), .ZN(n830) );
  NAND2_X1 U713 ( .A1(DATA1[20]), .A2(net76065), .ZN(n831) );
  OAI21_X1 U714 ( .B1(net76493), .B2(DATA2[20]), .A(net76161), .ZN(n828) );
  OAI21_X1 U715 ( .B1(n1630), .B2(n522), .A(n832), .ZN(n825) );
  AOI22_X1 U716 ( .A1(n661), .A2(n1569), .B1(net74123), .B2(n639), .ZN(n832)
         );
  NOR2_X1 U717 ( .A1(n833), .A2(n754), .ZN(n486) );
  NOR2_X1 U718 ( .A1(net74118), .A2(net74263), .ZN(n754) );
  NOR2_X1 U719 ( .A1(n834), .A2(n835), .ZN(n823) );
  OAI21_X1 U720 ( .B1(net74162), .B2(n1606), .A(n836), .ZN(n835) );
  AOI22_X1 U721 ( .A1(net74095), .A2(n1442), .B1(N1630), .B2(net76177), .ZN(
        n836) );
  OAI21_X1 U722 ( .B1(n496), .B2(net74128), .A(n837), .ZN(n834) );
  AOI22_X1 U723 ( .A1(net76479), .A2(n635), .B1(n514), .B2(n642), .ZN(n837) );
  AOI21_X1 U724 ( .B1(n563), .B2(n519), .A(n833), .ZN(n496) );
  OAI21_X1 U725 ( .B1(n1589), .B2(n1695), .A(n838), .ZN(n833) );
  AOI22_X1 U726 ( .A1(n1511), .A2(n839), .B1(net76542), .B2(n374), .ZN(n838)
         );
  AOI22_X1 U727 ( .A1(n263), .A2(net76163), .B1(net76554), .B2(n265), .ZN(n840) );
  NAND2_X1 U728 ( .A1(n841), .A2(n842), .ZN(n263) );
  NOR4_X1 U729 ( .A1(n843), .A2(n844), .A3(n845), .A4(n846), .ZN(n842) );
  AOI21_X1 U730 ( .B1(n847), .B2(net76161), .A(n1671), .ZN(n846) );
  AOI22_X1 U731 ( .A1(DATA1[19]), .A2(net76063), .B1(net76147), .B2(n1611), 
        .ZN(n847) );
  NOR2_X1 U732 ( .A1(n1653), .A2(n1685), .ZN(n845) );
  OAI21_X1 U733 ( .B1(n848), .B2(n1611), .A(net74292), .ZN(n844) );
  AOI21_X1 U734 ( .B1(net76149), .B2(n1671), .A(net76488), .ZN(n848) );
  OAI21_X1 U735 ( .B1(n1632), .B2(n522), .A(n849), .ZN(n843) );
  AOI22_X1 U736 ( .A1(n661), .A2(n1577), .B1(net74123), .B2(n398), .ZN(n849)
         );
  AOI21_X1 U737 ( .B1(n1578), .B2(n563), .A(n850), .ZN(n547) );
  NOR2_X1 U738 ( .A1(n851), .A2(n852), .ZN(n841) );
  OAI21_X1 U739 ( .B1(net74162), .B2(n1610), .A(n853), .ZN(n852) );
  AOI22_X1 U740 ( .A1(net74095), .A2(n1439), .B1(N1629), .B2(net76177), .ZN(
        n853) );
  OAI21_X1 U741 ( .B1(n564), .B2(net74128), .A(n854), .ZN(n851) );
  AOI22_X1 U742 ( .A1(net76479), .A2(n666), .B1(net76501), .B2(n524), .ZN(n854) );
  NAND2_X1 U743 ( .A1(n855), .A2(n856), .ZN(n524) );
  AOI22_X1 U744 ( .A1(DATA1[18]), .A2(net76067), .B1(DATA1[19]), .B2(n1527), 
        .ZN(n856) );
  AOI22_X1 U745 ( .A1(DATA1[16]), .A2(net76087), .B1(DATA1[17]), .B2(net76781), 
        .ZN(n855) );
  OAI21_X1 U747 ( .B1(net74244), .B2(n1693), .A(n857), .ZN(n850) );
  AOI22_X1 U748 ( .A1(net76542), .A2(n409), .B1(n465), .B2(n753), .ZN(n857) );
  AOI22_X1 U749 ( .A1(n265), .A2(net76163), .B1(net76555), .B2(n266), .ZN(n858) );
  NAND2_X1 U750 ( .A1(n859), .A2(n860), .ZN(n265) );
  NOR4_X1 U751 ( .A1(n861), .A2(n862), .A3(n863), .A4(n864), .ZN(n860) );
  AOI21_X1 U752 ( .B1(n865), .B2(net76161), .A(n1672), .ZN(n864) );
  AOI22_X1 U753 ( .A1(DATA1[18]), .A2(net76063), .B1(net76147), .B2(n1614), 
        .ZN(n865) );
  NOR2_X1 U754 ( .A1(n1654), .A2(n1685), .ZN(n863) );
  OAI21_X1 U755 ( .B1(n866), .B2(n1614), .A(net74292), .ZN(n862) );
  AOI21_X1 U756 ( .B1(net76149), .B2(n1672), .A(net76488), .ZN(n866) );
  OAI21_X1 U757 ( .B1(n1634), .B2(n522), .A(n867), .ZN(n861) );
  AOI22_X1 U758 ( .A1(n661), .A2(n1568), .B1(net74123), .B2(n428), .ZN(n867)
         );
  AOI21_X1 U759 ( .B1(n577), .B2(n563), .A(n868), .ZN(n808) );
  NOR2_X1 U760 ( .A1(n869), .A2(n870), .ZN(n859) );
  OAI21_X1 U761 ( .B1(net74162), .B2(n1613), .A(n871), .ZN(n870) );
  AOI22_X1 U762 ( .A1(net74095), .A2(DATA2[2]), .B1(N1628), .B2(net76177), 
        .ZN(n871) );
  OAI21_X1 U763 ( .B1(n819), .B2(net74128), .A(n872), .ZN(n869) );
  AOI22_X1 U764 ( .A1(net76479), .A2(n688), .B1(n514), .B2(n593), .ZN(n872) );
  NAND2_X1 U765 ( .A1(n873), .A2(n874), .ZN(n593) );
  AOI22_X1 U766 ( .A1(DATA1[17]), .A2(net76067), .B1(DATA1[18]), .B2(n1528), 
        .ZN(n874) );
  AOI22_X1 U767 ( .A1(DATA1[15]), .A2(net76089), .B1(DATA1[16]), .B2(net76778), 
        .ZN(n873) );
  AOI21_X1 U768 ( .B1(n578), .B2(net76535), .A(n868), .ZN(n819) );
  OAI21_X1 U769 ( .B1(n1585), .B2(n1693), .A(n875), .ZN(n868) );
  AOI22_X1 U770 ( .A1(net76542), .A2(n438), .B1(n465), .B2(n776), .ZN(n875) );
  AOI22_X1 U771 ( .A1(n266), .A2(net76163), .B1(net76554), .B2(n267), .ZN(n876) );
  NAND2_X1 U772 ( .A1(n877), .A2(n878), .ZN(n266) );
  NOR4_X1 U773 ( .A1(n879), .A2(n880), .A3(n881), .A4(n882), .ZN(n878) );
  AOI21_X1 U774 ( .B1(n883), .B2(net76161), .A(n1674), .ZN(n882) );
  AOI22_X1 U775 ( .A1(DATA1[17]), .A2(net76063), .B1(net76147), .B2(n1617), 
        .ZN(n883) );
  AOI21_X1 U776 ( .B1(n884), .B2(n885), .A(n627), .ZN(n881) );
  AOI22_X1 U777 ( .A1(net76542), .A2(n335), .B1(n465), .B2(n336), .ZN(n884) );
  NOR2_X1 U778 ( .A1(n1648), .A2(n747), .ZN(n880) );
  OAI21_X1 U779 ( .B1(n462), .B2(n1685), .A(n886), .ZN(n879) );
  AOI21_X1 U780 ( .B1(DATA1[17]), .B2(n887), .A(n650), .ZN(n886) );
  OAI21_X1 U781 ( .B1(DATA2[17]), .B2(net76493), .A(net76161), .ZN(n887) );
  NOR2_X1 U782 ( .A1(n888), .A2(n889), .ZN(n877) );
  OAI21_X1 U783 ( .B1(net74162), .B2(n1616), .A(n890), .ZN(n889) );
  AOI22_X1 U784 ( .A1(net74095), .A2(n1420), .B1(N1627), .B2(net76177), .ZN(
        n890) );
  OAI21_X1 U785 ( .B1(n1618), .B2(net74121), .A(n891), .ZN(n888) );
  AOI22_X1 U786 ( .A1(net74124), .A2(n346), .B1(n512), .B2(n611), .ZN(n891) );
  NAND2_X1 U787 ( .A1(n892), .A2(n893), .ZN(n610) );
  AOI22_X1 U788 ( .A1(DATA1[16]), .A2(net76071), .B1(DATA1[17]), .B2(n1528), 
        .ZN(n893) );
  AOI22_X1 U789 ( .A1(DATA1[14]), .A2(net76087), .B1(DATA1[15]), .B2(net76781), 
        .ZN(n892) );
  OAI21_X1 U790 ( .B1(n894), .B2(net76167), .A(n895), .ZN(OUTALU[15]) );
  NAND2_X1 U791 ( .A1(n267), .A2(net76165), .ZN(n895) );
  NAND2_X1 U792 ( .A1(n896), .A2(n897), .ZN(n267) );
  NOR4_X1 U793 ( .A1(n898), .A2(n899), .A3(n900), .A4(n901), .ZN(n897) );
  AOI22_X1 U795 ( .A1(DATA1[16]), .A2(net76065), .B1(net76147), .B2(n1621), 
        .ZN(n902) );
  AOI21_X1 U796 ( .B1(n903), .B2(n1582), .A(n627), .ZN(n900) );
  NOR2_X1 U797 ( .A1(n661), .A2(n703), .ZN(n627) );
  NOR2_X1 U798 ( .A1(n1701), .A2(n1442), .ZN(n703) );
  NOR2_X1 U799 ( .A1(n904), .A2(net74101), .ZN(n661) );
  AOI22_X1 U800 ( .A1(net76542), .A2(n381), .B1(n465), .B2(n374), .ZN(n903) );
  NOR2_X1 U801 ( .A1(n1650), .A2(n747), .ZN(n899) );
  NAND2_X1 U802 ( .A1(n1517), .A2(n582), .ZN(n747) );
  NAND2_X1 U803 ( .A1(n906), .A2(n907), .ZN(n898) );
  AOI21_X1 U804 ( .B1(n908), .B2(n519), .A(n650), .ZN(n907) );
  NOR2_X1 U805 ( .A1(n909), .A2(net74101), .ZN(n650) );
  NOR2_X1 U806 ( .A1(n1701), .A2(net74133), .ZN(n908) );
  AOI22_X1 U807 ( .A1(DATA1[16]), .A2(n910), .B1(n658), .B2(n723), .ZN(n906)
         );
  NOR2_X1 U808 ( .A1(net74133), .A2(n1700), .ZN(n658) );
  OAI21_X1 U809 ( .B1(DATA2[16]), .B2(net76493), .A(net76161), .ZN(n910) );
  NOR2_X1 U810 ( .A1(n911), .A2(n912), .ZN(n896) );
  OAI21_X1 U811 ( .B1(net74162), .B2(n1620), .A(n913), .ZN(n912) );
  AOI22_X1 U812 ( .A1(net74095), .A2(n1416), .B1(N1626), .B2(net76177), .ZN(
        n913) );
  OAI21_X1 U813 ( .B1(n1623), .B2(net74121), .A(n914), .ZN(n911) );
  AOI22_X1 U814 ( .A1(net74124), .A2(n639), .B1(n512), .B2(n636), .ZN(n914) );
  NOR2_X1 U815 ( .A1(n1692), .A2(n1700), .ZN(n512) );
  NAND2_X1 U816 ( .A1(n1520), .A2(n582), .ZN(n522) );
  OAI21_X1 U817 ( .B1(n915), .B2(net76169), .A(n916), .ZN(OUTALU[14]) );
  NOR4_X1 U819 ( .A1(n917), .A2(n918), .A3(n919), .A4(n920), .ZN(n894) );
  AOI21_X1 U820 ( .B1(n921), .B2(net76161), .A(net74147), .ZN(n920) );
  AOI22_X1 U821 ( .A1(DATA1[15]), .A2(net76065), .B1(net76147), .B2(n1624), 
        .ZN(n921) );
  AOI21_X1 U822 ( .B1(n922), .B2(n923), .A(n1701), .ZN(n919) );
  AOI21_X1 U823 ( .B1(n361), .B2(n409), .A(n924), .ZN(n923) );
  OAI21_X1 U824 ( .B1(n1619), .B2(net74119), .A(n925), .ZN(n924) );
  AOI22_X1 U826 ( .A1(n1520), .A2(n753), .B1(n1517), .B2(n926), .ZN(n922) );
  OAI21_X1 U827 ( .B1(n927), .B2(n1624), .A(n1571), .ZN(n918) );
  AOI21_X1 U828 ( .B1(net76149), .B2(net74147), .A(net76488), .ZN(n927) );
  NAND2_X1 U829 ( .A1(n928), .A2(n929), .ZN(n917) );
  AOI22_X1 U830 ( .A1(n411), .A2(n930), .B1(n535), .B2(n1434), .ZN(n929) );
  NAND2_X1 U831 ( .A1(n931), .A2(n932), .ZN(n535) );
  AOI22_X1 U832 ( .A1(net76542), .A2(n666), .B1(n563), .B2(n566), .ZN(n932) );
  NAND2_X1 U833 ( .A1(n933), .A2(n934), .ZN(n666) );
  AOI22_X1 U834 ( .A1(DATA1[14]), .A2(net76069), .B1(DATA1[15]), .B2(n1528), 
        .ZN(n934) );
  AOI22_X1 U835 ( .A1(DATA1[12]), .A2(net76087), .B1(DATA1[13]), .B2(net76778), 
        .ZN(n933) );
  AOI22_X1 U836 ( .A1(n1511), .A2(n398), .B1(n465), .B2(n659), .ZN(n931) );
  OR2_X1 U837 ( .A1(n935), .A2(n936), .ZN(n930) );
  NAND2_X1 U838 ( .A1(n937), .A2(n938), .ZN(n936) );
  AOI22_X1 U839 ( .A1(n1680), .A2(n753), .B1(n1681), .B2(n926), .ZN(n937) );
  OAI21_X1 U840 ( .B1(n1619), .B2(n333), .A(n939), .ZN(n935) );
  AOI22_X1 U841 ( .A1(n940), .A2(n1578), .B1(n1682), .B2(n409), .ZN(n939) );
  AOI22_X1 U842 ( .A1(N1625), .A2(net76177), .B1(N1994), .B2(net76506), .ZN(
        n928) );
  OAI21_X1 U843 ( .B1(n941), .B2(net76169), .A(n942), .ZN(OUTALU[13]) );
  NOR4_X1 U845 ( .A1(n943), .A2(n944), .A3(n945), .A4(n946), .ZN(n915) );
  AOI21_X1 U846 ( .B1(n947), .B2(net76161), .A(n1675), .ZN(n946) );
  AOI22_X1 U847 ( .A1(DATA1[14]), .A2(net76065), .B1(net76147), .B2(n1625), 
        .ZN(n947) );
  AOI21_X1 U848 ( .B1(n948), .B2(n949), .A(n1701), .ZN(n945) );
  AOI21_X1 U849 ( .B1(n361), .B2(n438), .A(n950), .ZN(n949) );
  OAI21_X1 U850 ( .B1(n1566), .B2(net74133), .A(n951), .ZN(n950) );
  NAND2_X1 U851 ( .A1(n405), .A2(n437), .ZN(n951) );
  AOI22_X1 U852 ( .A1(n1520), .A2(n776), .B1(n1517), .B2(n774), .ZN(n948) );
  OAI21_X1 U853 ( .B1(n952), .B2(n1625), .A(n1571), .ZN(n944) );
  AOI21_X1 U854 ( .B1(net76149), .B2(n1675), .A(net76487), .ZN(n952) );
  NAND2_X1 U855 ( .A1(n953), .A2(n954), .ZN(n943) );
  AOI22_X1 U856 ( .A1(n411), .A2(n955), .B1(n594), .B2(n1434), .ZN(n954) );
  NAND2_X1 U857 ( .A1(n956), .A2(n957), .ZN(n594) );
  AOI22_X1 U858 ( .A1(net76542), .A2(n688), .B1(n563), .B2(n781), .ZN(n957) );
  NAND2_X1 U859 ( .A1(n958), .A2(n959), .ZN(n688) );
  AOI21_X1 U860 ( .B1(DATA1[13]), .B2(net76069), .A(n960), .ZN(n959) );
  AOI22_X1 U861 ( .A1(DATA1[14]), .A2(n1527), .B1(DATA1[11]), .B2(net76087), 
        .ZN(n958) );
  AOI22_X1 U862 ( .A1(n1511), .A2(n428), .B1(n465), .B2(n682), .ZN(n956) );
  OR2_X1 U863 ( .A1(n961), .A2(n962), .ZN(n955) );
  NAND2_X1 U864 ( .A1(n963), .A2(n938), .ZN(n962) );
  AOI22_X1 U865 ( .A1(n1680), .A2(n776), .B1(n1681), .B2(n774), .ZN(n963) );
  OAI21_X1 U866 ( .B1(n1609), .B2(n964), .A(n965), .ZN(n961) );
  AOI22_X1 U867 ( .A1(n940), .A2(n577), .B1(n1679), .B2(n437), .ZN(n965) );
  AOI22_X1 U868 ( .A1(N1624), .A2(net76177), .B1(N1993), .B2(net76505), .ZN(
        n953) );
  OAI21_X1 U869 ( .B1(n966), .B2(net76169), .A(n967), .ZN(OUTALU[12]) );
  NAND2_X1 U870 ( .A1(n1559), .A2(net76167), .ZN(n967) );
  NOR4_X1 U871 ( .A1(n968), .A2(n1572), .A3(n969), .A4(n970), .ZN(n941) );
  AOI21_X1 U872 ( .B1(n971), .B2(n972), .A(n1701), .ZN(n970) );
  AOI21_X1 U873 ( .B1(n1517), .B2(n460), .A(n973), .ZN(n972) );
  OAI21_X1 U874 ( .B1(n1576), .B2(net74133), .A(n974), .ZN(n973) );
  NAND2_X1 U875 ( .A1(n405), .A2(n337), .ZN(n974) );
  AOI22_X1 U876 ( .A1(n361), .A2(n335), .B1(n1520), .B2(n336), .ZN(n971) );
  AOI21_X1 U877 ( .B1(n975), .B2(n1647), .A(n1690), .ZN(n969) );
  OAI21_X1 U878 ( .B1(n1648), .B2(n1693), .A(n976), .ZN(n614) );
  NAND2_X1 U879 ( .A1(n563), .A2(n1656), .ZN(n976) );
  NAND2_X1 U880 ( .A1(n977), .A2(n978), .ZN(n800) );
  AOI22_X1 U881 ( .A1(n1449), .A2(net76069), .B1(DATA1[5]), .B2(n1528), .ZN(
        n978) );
  AOI22_X1 U882 ( .A1(n1446), .A2(net76087), .B1(n1448), .B2(net76781), .ZN(
        n977) );
  AOI22_X1 U883 ( .A1(net76542), .A2(n611), .B1(n465), .B2(n346), .ZN(n975) );
  NAND2_X1 U884 ( .A1(n979), .A2(n980), .ZN(n346) );
  AOI22_X1 U885 ( .A1(DATA1[8]), .A2(net76069), .B1(DATA1[9]), .B2(n1528), 
        .ZN(n980) );
  AOI22_X1 U886 ( .A1(DATA1[6]), .A2(net76087), .B1(DATA1[7]), .B2(net76778), 
        .ZN(n979) );
  NAND2_X1 U887 ( .A1(n981), .A2(n982), .ZN(n611) );
  AOI22_X1 U888 ( .A1(DATA1[12]), .A2(net76069), .B1(DATA1[13]), .B2(n1528), 
        .ZN(n982) );
  AOI22_X1 U889 ( .A1(DATA1[10]), .A2(net76087), .B1(DATA1[11]), .B2(net76781), 
        .ZN(n981) );
  AOI21_X1 U890 ( .B1(n984), .B2(DATA1[13]), .A(n344), .ZN(n983) );
  OAI21_X1 U891 ( .B1(net76493), .B2(n1428), .A(net76161), .ZN(n984) );
  NAND2_X1 U892 ( .A1(n985), .A2(n986), .ZN(n968) );
  AOI22_X1 U893 ( .A1(n1428), .A2(n987), .B1(n411), .B2(n988), .ZN(n986) );
  OR2_X1 U894 ( .A1(n989), .A2(n990), .ZN(n988) );
  NAND2_X1 U895 ( .A1(n991), .A2(n938), .ZN(n990) );
  AOI22_X1 U896 ( .A1(n1681), .A2(n460), .B1(n1679), .B2(n337), .ZN(n991) );
  OAI21_X1 U897 ( .B1(n1597), .B2(n492), .A(n992), .ZN(n989) );
  AOI22_X1 U898 ( .A1(n940), .A2(n360), .B1(n1682), .B2(n335), .ZN(n992) );
  NAND2_X1 U899 ( .A1(n993), .A2(net76161), .ZN(n987) );
  AOI22_X1 U900 ( .A1(DATA1[13]), .A2(net76065), .B1(net76147), .B2(n1627), 
        .ZN(n993) );
  AOI22_X1 U901 ( .A1(N1623), .A2(net76177), .B1(N1992), .B2(net76507), .ZN(
        n985) );
  OAI21_X1 U902 ( .B1(n292), .B2(net76171), .A(n994), .ZN(OUTALU[11]) );
  NAND2_X1 U903 ( .A1(n1539), .A2(net76167), .ZN(n994) );
  NOR4_X1 U904 ( .A1(n995), .A2(n996), .A3(n997), .A4(n1558), .ZN(n966) );
  OAI21_X1 U905 ( .B1(n999), .B2(n1000), .A(n411), .ZN(n998) );
  NAND2_X1 U906 ( .A1(n1001), .A2(n938), .ZN(n1000) );
  AOI21_X1 U907 ( .B1(n445), .B2(n1002), .A(n418), .ZN(n938) );
  NOR2_X1 U908 ( .A1(net74263), .A2(net76542), .ZN(n1002) );
  AOI22_X1 U909 ( .A1(n1681), .A2(n735), .B1(n1679), .B2(n491), .ZN(n1001) );
  OAI21_X1 U910 ( .B1(n1602), .B2(n492), .A(n1003), .ZN(n999) );
  AOI22_X1 U911 ( .A1(n940), .A2(n839), .B1(n1682), .B2(n381), .ZN(n1003) );
  NOR2_X1 U912 ( .A1(n1683), .A2(net74115), .ZN(n940) );
  AOI21_X1 U913 ( .B1(n1004), .B2(net76161), .A(n1676), .ZN(n997) );
  AOI22_X1 U914 ( .A1(DATA1[12]), .A2(net76065), .B1(net76147), .B2(n1629), 
        .ZN(n1004) );
  OAI21_X1 U915 ( .B1(n1005), .B2(n1629), .A(n1571), .ZN(n996) );
  AOI21_X1 U916 ( .B1(net76149), .B2(n1676), .A(net76487), .ZN(n1005) );
  NAND2_X1 U917 ( .A1(n1006), .A2(n1007), .ZN(n995) );
  AOI22_X1 U918 ( .A1(n1008), .A2(n1434), .B1(n1009), .B2(n350), .ZN(n1007) );
  OR2_X1 U919 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
  OAI21_X1 U920 ( .B1(n1615), .B2(n1692), .A(n1012), .ZN(n1011) );
  AOI22_X1 U921 ( .A1(n1517), .A2(n735), .B1(n1520), .B2(n374), .ZN(n1012) );
  OAI21_X1 U922 ( .B1(n1626), .B2(net74119), .A(n1013), .ZN(n1010) );
  AOI22_X1 U923 ( .A1(n519), .A2(n359), .B1(n456), .B2(n839), .ZN(n1013) );
  OAI21_X1 U924 ( .B1(n1640), .B2(n1695), .A(n1014), .ZN(n1008) );
  AOI22_X1 U925 ( .A1(n1649), .A2(n1439), .B1(net76542), .B2(n636), .ZN(n1014)
         );
  OAI21_X1 U926 ( .B1(n723), .B2(n1696), .A(n1015), .ZN(n485) );
  NAND2_X1 U927 ( .A1(n1650), .A2(n1696), .ZN(n1015) );
  AOI22_X1 U928 ( .A1(N1622), .A2(net76177), .B1(N1991), .B2(net76506), .ZN(
        n1006) );
  OAI21_X1 U929 ( .B1(net76553), .B2(n292), .A(n1016), .ZN(OUTALU[10]) );
  NAND2_X1 U930 ( .A1(net76555), .A2(n291), .ZN(n1016) );
  OAI21_X1 U933 ( .B1(n1426), .B2(net76493), .A(net76161), .ZN(n1022) );
  NAND2_X1 U934 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
  OAI21_X1 U935 ( .B1(n1025), .B2(n1026), .A(n1027), .ZN(n1024) );
  OAI21_X1 U936 ( .B1(n684), .B2(n1683), .A(n1028), .ZN(n1026) );
  AOI22_X1 U937 ( .A1(n1680), .A2(n438), .B1(n1681), .B2(n776), .ZN(n1028) );
  AOI21_X1 U938 ( .B1(n577), .B2(n1509), .A(n1563), .ZN(n684) );
  AOI21_X1 U939 ( .B1(net76542), .B2(n774), .A(n707), .ZN(n1029) );
  OAI21_X1 U940 ( .B1(net74263), .B2(n1697), .A(n1030), .ZN(n577) );
  OAI21_X1 U941 ( .B1(n1622), .B2(n964), .A(n1031), .ZN(n1025) );
  AOI21_X1 U942 ( .B1(n1679), .B2(n432), .A(n418), .ZN(n1031) );
  AOI22_X1 U943 ( .A1(n397), .A2(n682), .B1(n1426), .B2(n1032), .ZN(n1019) );
  NAND2_X1 U944 ( .A1(n1033), .A2(net76161), .ZN(n1032) );
  AOI22_X1 U945 ( .A1(DATA1[10]), .A2(net76065), .B1(net76147), .B2(net74191), 
        .ZN(n1033) );
  NAND2_X1 U946 ( .A1(n1034), .A2(n1035), .ZN(n682) );
  AOI22_X1 U947 ( .A1(DATA1[9]), .A2(net76069), .B1(DATA1[10]), .B2(n1528), 
        .ZN(n1035) );
  AOI22_X1 U948 ( .A1(DATA1[7]), .A2(net76087), .B1(DATA1[8]), .B2(net76778), 
        .ZN(n1034) );
  AOI22_X1 U949 ( .A1(n681), .A2(n1434), .B1(n1036), .B2(n350), .ZN(n1018) );
  OR2_X1 U950 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
  OAI21_X1 U951 ( .B1(n1585), .B2(net74133), .A(n1039), .ZN(n1038) );
  AOI22_X1 U952 ( .A1(n1520), .A2(n438), .B1(n1517), .B2(n776), .ZN(n1039) );
  NAND2_X1 U953 ( .A1(n1040), .A2(n1041), .ZN(n776) );
  AOI22_X1 U954 ( .A1(DATA1[22]), .A2(net76069), .B1(DATA1[21]), .B2(n1528), 
        .ZN(n1041) );
  AOI22_X1 U955 ( .A1(DATA1[24]), .A2(net76087), .B1(DATA1[23]), .B2(net76781), 
        .ZN(n1040) );
  NAND2_X1 U956 ( .A1(n1042), .A2(n1043), .ZN(n438) );
  AOI22_X1 U957 ( .A1(DATA1[18]), .A2(net76069), .B1(DATA1[17]), .B2(n1528), 
        .ZN(n1043) );
  AOI22_X1 U958 ( .A1(DATA1[20]), .A2(net76087), .B1(DATA1[19]), .B2(net76778), 
        .ZN(n1042) );
  NAND2_X1 U959 ( .A1(n1044), .A2(n1045), .ZN(n774) );
  AOI22_X1 U960 ( .A1(DATA1[26]), .A2(net76069), .B1(DATA1[25]), .B2(n1527), 
        .ZN(n1045) );
  AOI22_X1 U961 ( .A1(net76087), .A2(DATA1[28]), .B1(DATA1[27]), .B2(net76781), 
        .ZN(n1044) );
  OAI21_X1 U962 ( .B1(n1622), .B2(n1692), .A(n1046), .ZN(n1037) );
  AOI22_X1 U963 ( .A1(n359), .A2(n578), .B1(n405), .B2(n432), .ZN(n1046) );
  NAND2_X1 U964 ( .A1(n1047), .A2(n1048), .ZN(n432) );
  AOI22_X1 U965 ( .A1(DATA1[10]), .A2(net76069), .B1(DATA1[9]), .B2(n1527), 
        .ZN(n1048) );
  AOI22_X1 U966 ( .A1(DATA1[12]), .A2(net76087), .B1(DATA1[11]), .B2(net76107), 
        .ZN(n1047) );
  OAI21_X1 U967 ( .B1(net74263), .B2(net81902), .A(n1030), .ZN(n578) );
  NOR2_X1 U969 ( .A1(n1435), .A2(net74246), .ZN(n1049) );
  NAND2_X1 U970 ( .A1(n1050), .A2(n1051), .ZN(n437) );
  AOI22_X1 U971 ( .A1(DATA1[14]), .A2(net76069), .B1(DATA1[13]), .B2(n1527), 
        .ZN(n1051) );
  AOI22_X1 U972 ( .A1(DATA1[16]), .A2(net76087), .B1(DATA1[15]), .B2(net76107), 
        .ZN(n1050) );
  OAI21_X1 U973 ( .B1(n1644), .B2(n1695), .A(n1052), .ZN(n681) );
  NAND2_X1 U974 ( .A1(n562), .A2(n781), .ZN(n1052) );
  OAI21_X1 U975 ( .B1(net81902), .B2(n1660), .A(n1053), .ZN(n781) );
  NOR2_X1 U976 ( .A1(n1054), .A2(n555), .ZN(n1053) );
  NOR2_X1 U977 ( .A1(n1655), .A2(n1435), .ZN(n555) );
  NAND2_X1 U978 ( .A1(n1055), .A2(n1056), .ZN(n428) );
  AOI21_X1 U979 ( .B1(DATA1[5]), .B2(net76069), .A(n1057), .ZN(n1056) );
  AOI21_X1 U980 ( .B1(DATA1[6]), .B2(n1527), .A(n557), .ZN(n1055) );
  NOR2_X1 U981 ( .A1(n1651), .A2(net81902), .ZN(n557) );
  AOI22_X1 U982 ( .A1(N1620), .A2(net76177), .B1(N1989), .B2(net76505), .ZN(
        n1017) );
  NOR4_X1 U983 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n292) );
  AOI21_X1 U984 ( .B1(n1062), .B2(n1557), .A(n1662), .ZN(n1061) );
  NOR2_X1 U985 ( .A1(n1663), .A2(net74101), .ZN(n411) );
  OAI21_X1 U986 ( .B1(n964), .B2(n1619), .A(n1064), .ZN(n1063) );
  AOI21_X1 U987 ( .B1(n402), .B2(n1679), .A(n418), .ZN(n1064) );
  NAND2_X1 U988 ( .A1(n1065), .A2(n1509), .ZN(n964) );
  AOI21_X1 U989 ( .B1(n445), .B2(n662), .A(n1066), .ZN(n1062) );
  OAI21_X1 U990 ( .B1(n1605), .B2(n492), .A(n1067), .ZN(n1066) );
  NAND2_X1 U991 ( .A1(n1681), .A2(n753), .ZN(n1067) );
  NAND2_X1 U992 ( .A1(n1065), .A2(n563), .ZN(n415) );
  NAND2_X1 U993 ( .A1(n1065), .A2(n562), .ZN(n492) );
  OAI21_X1 U994 ( .B1(n1068), .B2(n1695), .A(n1069), .ZN(n662) );
  AOI21_X1 U995 ( .B1(net76542), .B2(n926), .A(n707), .ZN(n1069) );
  NOR2_X1 U996 ( .A1(n1694), .A2(net74263), .ZN(n707) );
  NOR2_X1 U997 ( .A1(n1684), .A2(n1687), .ZN(n445) );
  AOI22_X1 U999 ( .A1(DATA1[11]), .A2(net76065), .B1(net76147), .B2(n1631), 
        .ZN(n1070) );
  OAI21_X1 U1000 ( .B1(n1632), .B2(n1689), .A(n1071), .ZN(n1059) );
  AOI21_X1 U1001 ( .B1(DATA1[11]), .B2(n1072), .A(n344), .ZN(n1071) );
  NOR2_X1 U1002 ( .A1(n1023), .A2(net74101), .ZN(n344) );
  AOI21_X1 U1003 ( .B1(n1073), .B2(net76578), .A(n1579), .ZN(n1023) );
  OAI21_X1 U1004 ( .B1(net82738), .B2(net76493), .A(net76159), .ZN(n1072) );
  NOR2_X1 U1005 ( .A1(net74115), .A2(n1690), .ZN(n397) );
  NAND2_X1 U1006 ( .A1(n1074), .A2(n1075), .ZN(n659) );
  AOI22_X1 U1007 ( .A1(DATA1[10]), .A2(net76069), .B1(DATA1[11]), .B2(n1527), 
        .ZN(n1075) );
  AOI22_X1 U1008 ( .A1(DATA1[8]), .A2(net76089), .B1(DATA1[9]), .B2(net76781), 
        .ZN(n1074) );
  NAND2_X1 U1009 ( .A1(n1076), .A2(n1077), .ZN(n1058) );
  AOI22_X1 U1010 ( .A1(n657), .A2(n1434), .B1(n1078), .B2(n350), .ZN(n1077) );
  OR2_X1 U1011 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
  OAI21_X1 U1012 ( .B1(net74244), .B2(net74133), .A(n1081), .ZN(n1080) );
  AOI22_X1 U1013 ( .A1(n1520), .A2(n409), .B1(n1517), .B2(n753), .ZN(n1081) );
  NAND2_X1 U1014 ( .A1(n1082), .A2(n1083), .ZN(n753) );
  AOI22_X1 U1015 ( .A1(DATA1[23]), .A2(net76071), .B1(DATA1[22]), .B2(n1527), 
        .ZN(n1083) );
  AOI22_X1 U1016 ( .A1(DATA1[25]), .A2(net76089), .B1(DATA1[24]), .B2(net76107), .ZN(n1082) );
  NAND2_X1 U1017 ( .A1(n1084), .A2(n1085), .ZN(n409) );
  AOI22_X1 U1018 ( .A1(DATA1[19]), .A2(net76071), .B1(DATA1[18]), .B2(n1530), 
        .ZN(n1085) );
  AOI22_X1 U1019 ( .A1(DATA1[21]), .A2(net76089), .B1(DATA1[20]), .B2(net76107), .ZN(n1084) );
  NAND2_X1 U1020 ( .A1(n1086), .A2(n1087), .ZN(n926) );
  AOI22_X1 U1021 ( .A1(DATA1[27]), .A2(net76071), .B1(DATA1[26]), .B2(n1530), 
        .ZN(n1087) );
  AOI22_X1 U1022 ( .A1(net76087), .A2(DATA1[29]), .B1(net76781), .B2(DATA1[28]), .ZN(n1086) );
  OAI21_X1 U1023 ( .B1(n1619), .B2(n1692), .A(n1088), .ZN(n1079) );
  NAND2_X1 U1025 ( .A1(n1089), .A2(n1090), .ZN(n402) );
  NOR2_X1 U1026 ( .A1(n1091), .A2(n960), .ZN(n1090) );
  NOR2_X1 U1027 ( .A1(n1629), .A2(net81902), .ZN(n960) );
  AOI22_X1 U1028 ( .A1(DATA1[11]), .A2(net76071), .B1(DATA1[10]), .B2(n1530), 
        .ZN(n1089) );
  AOI21_X1 U1029 ( .B1(net76578), .B2(net76069), .A(n591), .ZN(n652) );
  NAND2_X1 U1030 ( .A1(n1092), .A2(n1093), .ZN(n408) );
  AOI22_X1 U1031 ( .A1(DATA1[15]), .A2(net76071), .B1(DATA1[14]), .B2(n1527), 
        .ZN(n1093) );
  AOI22_X1 U1032 ( .A1(DATA1[17]), .A2(net76089), .B1(DATA1[16]), .B2(net76107), .ZN(n1092) );
  OAI33_X1 U1033 ( .A1(n1094), .A2(n1442), .A3(net83235), .B1(n1095), .B2(
        n1442), .B3(net83422), .ZN(n352) );
  OAI21_X1 U1034 ( .B1(n1653), .B2(n1693), .A(n1096), .ZN(n657) );
  NAND2_X1 U1035 ( .A1(n1509), .A2(n398), .ZN(n1096) );
  NAND2_X1 U1036 ( .A1(n1097), .A2(n1098), .ZN(n398) );
  AOI22_X1 U1037 ( .A1(DATA1[6]), .A2(net76071), .B1(DATA1[7]), .B2(n1530), 
        .ZN(n1098) );
  AOI22_X1 U1038 ( .A1(n1449), .A2(net76089), .B1(DATA1[5]), .B2(net76107), 
        .ZN(n1097) );
  NAND2_X1 U1039 ( .A1(n1099), .A2(n1100), .ZN(n566) );
  AOI22_X1 U1040 ( .A1(n1446), .A2(net76071), .B1(n1448), .B2(n1530), .ZN(
        n1100) );
  AOI22_X1 U1041 ( .A1(n1444), .A2(net76089), .B1(n1411), .B2(net76107), .ZN(
        n1099) );
  AOI22_X1 U1042 ( .A1(N1621), .A2(net76177), .B1(N1990), .B2(net76507), .ZN(
        n1076) );
  OAI21_X1 U1043 ( .B1(n289), .B2(net76171), .A(n1101), .ZN(OUTALU[0]) );
  NAND2_X1 U1044 ( .A1(n268), .A2(net76163), .ZN(n1101) );
  NAND2_X1 U1045 ( .A1(n1102), .A2(n1103), .ZN(n268) );
  NOR4_X1 U1046 ( .A1(n544), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1103) );
  AOI21_X1 U1047 ( .B1(n1107), .B2(net76161), .A(n1697), .ZN(n1106) );
  AOI22_X1 U1048 ( .A1(n1411), .A2(net76061), .B1(net76149), .B2(n1657), .ZN(
        n1107) );
  NOR2_X1 U1050 ( .A1(n1110), .A2(n1657), .ZN(n1105) );
  AOI21_X1 U1051 ( .B1(net76149), .B2(n1697), .A(net76487), .ZN(n1110) );
  OAI21_X1 U1052 ( .B1(net74096), .B2(n1094), .A(n1111), .ZN(net76487) );
  OR2_X1 U1053 ( .A1(n1109), .A2(net94830), .ZN(n1111) );
  NAND2_X1 U1054 ( .A1(n301), .A2(n1112), .ZN(n1109) );
  NAND2_X1 U1055 ( .A1(n301), .A2(n1113), .ZN(net76493) );
  OAI21_X1 U1056 ( .B1(net76573), .B2(n1114), .A(net74089), .ZN(n1113) );
  AOI21_X1 U1057 ( .B1(n1701), .B2(n546), .A(n1115), .ZN(n1104) );
  NOR4_X1 U1058 ( .A1(n1116), .A2(n1596), .A3(n1117), .A4(n1118), .ZN(n1115)
         );
  NOR2_X1 U1059 ( .A1(n1119), .A2(net74119), .ZN(n1118) );
  NOR4_X1 U1060 ( .A1(n1054), .A2(n723), .A3(n1057), .A4(n1120), .ZN(n1119) );
  NOR2_X1 U1061 ( .A1(net81902), .A2(n1655), .ZN(n1120) );
  NOR2_X1 U1062 ( .A1(n1652), .A2(n1704), .ZN(n1057) );
  NOR2_X1 U1063 ( .A1(n1657), .A2(n1703), .ZN(n1054) );
  NOR2_X1 U1064 ( .A1(n885), .A2(n1687), .ZN(n1117) );
  AOI21_X1 U1065 ( .B1(n360), .B2(net76535), .A(n1121), .ZN(n885) );
  NOR2_X1 U1066 ( .A1(n1693), .A2(n1587), .ZN(n1121) );
  NAND2_X1 U1067 ( .A1(n1122), .A2(n1123), .ZN(n460) );
  AOI22_X1 U1068 ( .A1(DATA1[25]), .A2(net76071), .B1(DATA1[24]), .B2(n1530), 
        .ZN(n1123) );
  AOI22_X1 U1069 ( .A1(DATA1[27]), .A2(net76089), .B1(DATA1[26]), .B2(net76107), .ZN(n1122) );
  NAND2_X1 U1070 ( .A1(n1124), .A2(n1125), .ZN(n360) );
  AOI22_X1 U1071 ( .A1(DATA1[29]), .A2(net76071), .B1(DATA1[28]), .B2(n1530), 
        .ZN(n1125) );
  AOI22_X1 U1072 ( .A1(net76087), .A2(net76578), .B1(DATA1[30]), .B2(net76107), 
        .ZN(n1124) );
  AOI21_X1 U1073 ( .B1(n337), .B2(n1517), .A(n1127), .ZN(n1126) );
  NOR2_X1 U1074 ( .A1(net74135), .A2(n1597), .ZN(n1127) );
  NAND2_X1 U1075 ( .A1(n1128), .A2(n1129), .ZN(n336) );
  AOI22_X1 U1076 ( .A1(DATA1[21]), .A2(net76069), .B1(DATA1[20]), .B2(n1530), 
        .ZN(n1129) );
  NOR2_X1 U1077 ( .A1(n691), .A2(n1130), .ZN(n1128) );
  NOR2_X1 U1078 ( .A1(n1599), .A2(n1704), .ZN(n691) );
  NAND2_X1 U1079 ( .A1(n1131), .A2(n1132), .ZN(n337) );
  AOI22_X1 U1080 ( .A1(DATA1[13]), .A2(net76069), .B1(DATA1[12]), .B2(n1530), 
        .ZN(n1132) );
  AOI22_X1 U1081 ( .A1(DATA1[15]), .A2(net76091), .B1(DATA1[14]), .B2(net76107), .ZN(n1131) );
  OAI21_X1 U1082 ( .B1(n1633), .B2(n1691), .A(n1133), .ZN(n1116) );
  AOI22_X1 U1083 ( .A1(n361), .A2(n461), .B1(n456), .B2(n335), .ZN(n1133) );
  NAND2_X1 U1084 ( .A1(n1134), .A2(n1135), .ZN(n335) );
  AOI22_X1 U1085 ( .A1(DATA1[17]), .A2(net76069), .B1(DATA1[16]), .B2(n1530), 
        .ZN(n1135) );
  AOI22_X1 U1086 ( .A1(DATA1[19]), .A2(net76089), .B1(DATA1[18]), .B2(net76107), .ZN(n1134) );
  NAND2_X1 U1087 ( .A1(n1136), .A2(n1137), .ZN(n461) );
  AOI21_X1 U1088 ( .B1(DATA1[5]), .B2(net76069), .A(n1138), .ZN(n1137) );
  AOI22_X1 U1089 ( .A1(DATA1[7]), .A2(net76091), .B1(DATA1[6]), .B2(net76107), 
        .ZN(n1136) );
  NAND2_X1 U1090 ( .A1(n1139), .A2(n1140), .ZN(n473) );
  AOI22_X1 U1091 ( .A1(DATA1[9]), .A2(net76071), .B1(DATA1[8]), .B2(n1530), 
        .ZN(n1140) );
  AOI22_X1 U1092 ( .A1(DATA1[11]), .A2(net76089), .B1(DATA1[10]), .B2(net76107), .ZN(n1139) );
  NAND2_X1 U1093 ( .A1(n1141), .A2(n1142), .ZN(n546) );
  NOR2_X1 U1094 ( .A1(net74101), .A2(n1713), .ZN(n1141) );
  OAI21_X1 U1095 ( .B1(net83235), .B2(net74089), .A(n1143), .ZN(n350) );
  NAND2_X1 U1096 ( .A1(n1144), .A2(n315), .ZN(n1143) );
  NOR2_X1 U1098 ( .A1(net74101), .A2(n1146), .ZN(n544) );
  NOR4_X1 U1099 ( .A1(n1581), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1146)
         );
  AOI21_X1 U1100 ( .B1(N1980), .B2(net76506), .A(n1150), .ZN(n1102) );
  OAI21_X1 U1101 ( .B1(n462), .B2(net74121), .A(n1151), .ZN(n1150) );
  NAND2_X1 U1102 ( .A1(N1611), .A2(net76177), .ZN(n1151) );
  NOR2_X1 U1103 ( .A1(net74119), .A2(n1700), .ZN(n514) );
  NOR2_X1 U1104 ( .A1(n1152), .A2(n818), .ZN(n462) );
  NOR2_X1 U1105 ( .A1(n1657), .A2(n1435), .ZN(n818) );
  AOI21_X1 U1107 ( .B1(n301), .B2(net84449), .A(n1699), .ZN(n526) );
  AOI21_X1 U1108 ( .B1(n1155), .B2(n1156), .A(n1157), .ZN(n1154) );
  OAI21_X1 U1123 ( .B1(net76566), .B2(net74299), .A(n1173), .ZN(n1163) );
  AOI21_X1 U1125 ( .B1(net84454), .B2(net77259), .A(net82584), .ZN(n1174) );
  OAI21_X1 U1127 ( .B1(net76542), .B2(net74263), .A(n909), .ZN(n1176) );
  NOR4_X1 U1128 ( .A1(n1579), .A2(n1147), .A3(n1177), .A4(n1148), .ZN(n909) );
  OAI21_X1 U1129 ( .B1(net74263), .B2(n1671), .A(n1178), .ZN(n1148) );
  AOI21_X1 U1130 ( .B1(n1179), .B2(n1687), .A(net74263), .ZN(n1177) );
  OAI21_X1 U1131 ( .B1(n1673), .B2(net74263), .A(n1555), .ZN(n1147) );
  NOR2_X1 U1132 ( .A1(net74263), .A2(n1180), .ZN(n418) );
  NAND2_X1 U1133 ( .A1(n576), .A2(n1578), .ZN(n1175) );
  AOI21_X1 U1134 ( .B1(n1435), .B2(net76578), .A(n591), .ZN(n1068) );
  NOR2_X1 U1135 ( .A1(net74249), .A2(n1435), .ZN(n591) );
  NAND2_X1 U1136 ( .A1(n1183), .A2(n1065), .ZN(n904) );
  NOR2_X1 U1137 ( .A1(n1181), .A2(n1713), .ZN(n1183) );
  OAI21_X1 U1144 ( .B1(net76553), .B2(n289), .A(n1193), .ZN(CARRY) );
  NAND2_X1 U1145 ( .A1(net82056), .A2(net76554), .ZN(n1193) );
  AOI21_X1 U1148 ( .B1(n1155), .B2(n1201), .A(n1157), .ZN(n1200) );
  OAI21_X1 U1152 ( .B1(net76573), .B2(net83605), .A(n1158), .ZN(n1201) );
  OR2_X1 U1156 ( .A1(n528), .A2(n1159), .ZN(n1204) );
  NOR2_X1 U1157 ( .A1(n1205), .A2(net84454), .ZN(n1159) );
  OR2_X1 U1158 ( .A1(net83443), .A2(n311), .ZN(n1205) );
  NAND2_X1 U1159 ( .A1(n1206), .A2(n313), .ZN(n528) );
  NOR2_X1 U1162 ( .A1(n1435), .A2(net74263), .ZN(n519) );
  NAND2_X1 U1164 ( .A1(n1209), .A2(n301), .ZN(n510) );
  NOR2_X1 U1166 ( .A1(net76759), .A2(n1114), .ZN(n1209) );
  OAI21_X1 U1167 ( .B1(net74101), .B2(net74263), .A(n1210), .ZN(n1195) );
  OAI21_X1 U1168 ( .B1(n1211), .B2(n1212), .A(n582), .ZN(n1210) );
  OAI21_X1 U1169 ( .B1(net83422), .B2(n1095), .A(n1213), .ZN(n582) );
  OR2_X1 U1170 ( .A1(n1094), .A2(net83235), .ZN(n1213) );
  NAND2_X1 U1171 ( .A1(n1214), .A2(n1112), .ZN(n1095) );
  NOR2_X1 U1172 ( .A1(n1191), .A2(net83443), .ZN(n1112) );
  NOR2_X1 U1173 ( .A1(net76566), .A2(net76573), .ZN(n1214) );
  OAI21_X1 U1174 ( .B1(n1594), .B2(n1691), .A(n1215), .ZN(n1212) );
  AOI22_X1 U1175 ( .A1(n1517), .A2(n642), .B1(n456), .B2(n635), .ZN(n1215) );
  NAND2_X1 U1176 ( .A1(n1216), .A2(n1217), .ZN(n635) );
  AOI21_X1 U1177 ( .B1(DATA1[15]), .B2(net76071), .A(n1091), .ZN(n1217) );
  NOR2_X1 U1178 ( .A1(n1627), .A2(n1704), .ZN(n1091) );
  AOI22_X1 U1179 ( .A1(DATA1[16]), .A2(n1527), .B1(DATA1[14]), .B2(net76107), 
        .ZN(n1216) );
  NAND2_X1 U1180 ( .A1(n1218), .A2(n1219), .ZN(n642) );
  AOI22_X1 U1181 ( .A1(DATA1[19]), .A2(net76071), .B1(DATA1[20]), .B2(n1530), 
        .ZN(n1219) );
  AOI22_X1 U1182 ( .A1(DATA1[17]), .A2(net76091), .B1(DATA1[18]), .B2(net76107), .ZN(n1218) );
  NAND2_X1 U1183 ( .A1(n1220), .A2(n1221), .ZN(n733) );
  AOI21_X1 U1184 ( .B1(DATA1[23]), .B2(net76071), .A(n1130), .ZN(n1221) );
  NOR2_X1 U1185 ( .A1(n1601), .A2(net81902), .ZN(n1130) );
  AOI22_X1 U1186 ( .A1(DATA1[24]), .A2(n1527), .B1(DATA1[21]), .B2(net76087), 
        .ZN(n1220) );
  NAND2_X1 U1187 ( .A1(n1222), .A2(n1223), .ZN(n1211) );
  AOI22_X1 U1188 ( .A1(n1442), .A2(n1224), .B1(n405), .B2(n1225), .ZN(n1223)
         );
  OAI21_X1 U1189 ( .B1(net81902), .B2(net74249), .A(n1226), .ZN(n1225) );
  AOI22_X1 U1190 ( .A1(net76069), .A2(net76578), .B1(net76087), .B2(DATA1[29]), 
        .ZN(n1226) );
  OAI21_X1 U1191 ( .B1(n1640), .B2(n1693), .A(n1227), .ZN(n1224) );
  NAND2_X1 U1192 ( .A1(n563), .A2(n725), .ZN(n1227) );
  NAND2_X1 U1193 ( .A1(n1228), .A2(n1229), .ZN(n725) );
  AOI21_X1 U1194 ( .B1(n1411), .B2(net76087), .A(n1138), .ZN(n1229) );
  NOR2_X1 U1195 ( .A1(n1651), .A2(n1435), .ZN(n1138) );
  AOI21_X1 U1196 ( .B1(n1446), .B2(net76781), .A(n556), .ZN(n1228) );
  NOR2_X1 U1197 ( .A1(n1652), .A2(n1703), .ZN(n556) );
  NAND2_X1 U1198 ( .A1(n1230), .A2(n1231), .ZN(n639) );
  AOI22_X1 U1199 ( .A1(DATA1[7]), .A2(net76071), .B1(DATA1[8]), .B2(n1530), 
        .ZN(n1231) );
  AOI22_X1 U1200 ( .A1(DATA1[5]), .A2(net76091), .B1(DATA1[6]), .B2(net76107), 
        .ZN(n1230) );
  AOI22_X1 U1201 ( .A1(n359), .A2(n636), .B1(n361), .B2(n641), .ZN(n1222) );
  NAND2_X1 U1202 ( .A1(n1232), .A2(n1233), .ZN(n641) );
  AOI22_X1 U1203 ( .A1(DATA1[27]), .A2(net76071), .B1(DATA1[28]), .B2(n1530), 
        .ZN(n1233) );
  AOI22_X1 U1204 ( .A1(DATA1[25]), .A2(net76091), .B1(DATA1[26]), .B2(net76107), .ZN(n1232) );
  NAND2_X1 U1205 ( .A1(n1234), .A2(n1235), .ZN(n636) );
  AOI22_X1 U1206 ( .A1(DATA1[11]), .A2(net76071), .B1(DATA1[12]), .B2(n1530), 
        .ZN(n1235) );
  AOI22_X1 U1207 ( .A1(DATA1[9]), .A2(net76091), .B1(DATA1[10]), .B2(net76107), 
        .ZN(n1234) );
  NOR2_X1 U1211 ( .A1(n1239), .A2(n1240), .ZN(n289) );
  OAI21_X1 U1212 ( .B1(n1241), .B2(net83235), .A(n1242), .ZN(n1240) );
  AOI22_X1 U1213 ( .A1(n1155), .A2(n1243), .B1(N1610), .B2(net76177), .ZN(
        n1242) );
  OR2_X1 U1216 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
  OAI21_X1 U1217 ( .B1(N1577), .B2(n1094), .A(n1247), .ZN(n1246) );
  AOI22_X1 U1218 ( .A1(N1576), .A2(net74087), .B1(n1145), .B2(n1535), .ZN(
        n1247) );
  OAI21_X1 U1219 ( .B1(n1536), .B2(n313), .A(n1248), .ZN(n1245) );
  AOI21_X1 U1220 ( .B1(N1979), .B2(n1249), .A(n1250), .ZN(n1248) );
  NOR3_X1 U1221 ( .A1(n1702), .A2(n1537), .A3(net84454), .ZN(n1250) );
  OAI21_X1 U1223 ( .B1(net83262), .B2(n251), .A(n1192), .ZN(n1158) );
  NAND2_X1 U1224 ( .A1(n1253), .A2(net83262), .ZN(n1192) );
  NAND2_X1 U1226 ( .A1(net83262), .A2(n320), .ZN(n1252) );
  NOR2_X1 U1227 ( .A1(net82584), .A2(net83422), .ZN(n1155) );
  NOR3_X1 U1228 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1241) );
  OAI33_X1 U1229 ( .A1(n1659), .A2(net74119), .A3(n1094), .B1(n1108), .B2(
        n1698), .B3(n1660), .ZN(n1256) );
  NAND2_X1 U1230 ( .A1(n251), .A2(n252), .ZN(n1108) );
  NAND2_X1 U1231 ( .A1(n1257), .A2(n310), .ZN(n1094) );
  AOI21_X1 U1232 ( .B1(n1206), .B2(n313), .A(n1658), .ZN(n1255) );
  NAND2_X1 U1233 ( .A1(n314), .A2(n252), .ZN(n313) );
  OAI21_X1 U1234 ( .B1(n1258), .B2(n1236), .A(n1259), .ZN(n1254) );
  NAND2_X1 U1235 ( .A1(n1145), .A2(n1260), .ZN(n1259) );
  NOR2_X1 U1236 ( .A1(n1702), .A2(net82724), .ZN(n1145) );
  NAND2_X1 U1238 ( .A1(n1257), .A2(n314), .ZN(n1236) );
  NOR2_X1 U1239 ( .A1(net83262), .A2(net76573), .ZN(n1257) );
  OAI21_X1 U1240 ( .B1(n1261), .B2(net84454), .A(n1262), .ZN(n1239) );
  NOR2_X1 U1245 ( .A1(n1268), .A2(net82584), .ZN(n1267) );
  AOI21_X1 U1246 ( .B1(n321), .B2(n1535), .A(n1269), .ZN(n1268) );
  OAI33_X1 U1247 ( .A1(n1535), .A2(net83443), .A3(net76759), .B1(n1536), .B2(
        net76573), .B3(net77259), .ZN(n1269) );
  NOR3_X1 U1248 ( .A1(n1270), .A2(net76566), .A3(n321), .ZN(n1266) );
  NOR2_X1 U1249 ( .A1(net83443), .A2(net76573), .ZN(n321) );
  AOI22_X1 U1250 ( .A1(N1979), .A2(net74079), .B1(net82953), .B2(n1536), .ZN(
        n1270) );
  AOI21_X1 U1252 ( .B1(n1271), .B2(n1272), .A(net84429), .ZN(n1263) );
  AOI22_X1 U1253 ( .A1(n310), .A2(n1273), .B1(n1274), .B2(net81160), .ZN(n1272) );
  OAI21_X1 U1254 ( .B1(net76573), .B2(n1275), .A(n1276), .ZN(n1273) );
  AOI22_X1 U1255 ( .A1(n251), .A2(n1251), .B1(n314), .B2(n1277), .ZN(n1271) );
  OAI21_X1 U1256 ( .B1(net76573), .B2(n1538), .A(n1278), .ZN(n1251) );
  NAND2_X1 U1257 ( .A1(N1573), .A2(net76573), .ZN(n1278) );
  AOI21_X1 U1258 ( .B1(n1279), .B2(n315), .A(n1280), .ZN(n1261) );
  AOI21_X1 U1259 ( .B1(n1281), .B2(n1282), .A(net84429), .ZN(n1280) );
  OAI21_X1 U1260 ( .B1(n1283), .B2(n251), .A(N1979), .ZN(n1282) );
  NOR3_X1 U1261 ( .A1(n311), .A2(net76566), .A3(net83443), .ZN(n1283) );
  XNOR2_X1 U1262 ( .A(net76573), .B(n1284), .ZN(n311) );
  NOR4_X1 U1263 ( .A1(DATA2[31]), .A2(n1435), .A3(n333), .A4(n1663), .ZN(n1284) );
  NOR2_X1 U1264 ( .A1(n1073), .A2(n1185), .ZN(n1027) );
  NOR3_X1 U1266 ( .A1(DATA2[19]), .A2(DATA2[21]), .A3(DATA2[20]), .ZN(n1288)
         );
  NOR3_X1 U1267 ( .A1(n1428), .A2(DATA2[18]), .A3(n1430), .ZN(n1287) );
  NOR3_X1 U1268 ( .A1(n1669), .A2(n1424), .A3(net82738), .ZN(n1286) );
  NOR3_X1 U1269 ( .A1(n1667), .A2(n1290), .A3(n1291), .ZN(n1285) );
  NOR4_X1 U1270 ( .A1(DATA2[28]), .A2(DATA2[27]), .A3(DATA2[26]), .A4(
        DATA2[25]), .ZN(n1179) );
  NAND2_X1 U1271 ( .A1(n1065), .A2(net76542), .ZN(n333) );
  NOR2_X1 U1272 ( .A1(n1684), .A2(n1442), .ZN(n1065) );
  OAI21_X1 U1273 ( .B1(n1292), .B2(n1293), .A(net76566), .ZN(n1281) );
  NOR2_X1 U1274 ( .A1(n1294), .A2(n1702), .ZN(n1293) );
  AOI22_X1 U1275 ( .A1(net76573), .A2(n1661), .B1(n1444), .B2(n1416), .ZN(
        n1294) );
  NOR2_X1 U1276 ( .A1(n1416), .A2(n1444), .ZN(n1275) );
  XNOR2_X1 U1278 ( .A(n1444), .B(n1416), .ZN(n1276) );
  AOI21_X1 U1280 ( .B1(n1295), .B2(n1296), .A(net76566), .ZN(n1279) );
  AOI21_X1 U1281 ( .B1(n1297), .B2(n314), .A(n1298), .ZN(n1296) );
  NOR2_X1 U1282 ( .A1(net76573), .A2(n1299), .ZN(n1298) );
  AOI21_X1 U1283 ( .B1(n314), .B2(n1260), .A(n1300), .ZN(n1299) );
  NOR3_X1 U1284 ( .A1(n1659), .A2(net74119), .A3(n1702), .ZN(n1300) );
  NOR2_X1 U1285 ( .A1(net82953), .A2(net83443), .ZN(n310) );
  NOR2_X1 U1286 ( .A1(n1660), .A2(n1435), .ZN(n723) );
  NOR2_X1 U1287 ( .A1(net77259), .A2(net82953), .ZN(n314) );
  NOR2_X1 U1288 ( .A1(n1258), .A2(net76759), .ZN(n1297) );
  NOR2_X1 U1289 ( .A1(n1301), .A2(n1149), .ZN(n1258) );
  NAND2_X1 U1290 ( .A1(n1302), .A2(n1182), .ZN(n1149) );
  NAND2_X1 U1291 ( .A1(net76578), .A2(n1185), .ZN(n1182) );
  OAI21_X1 U1292 ( .B1(DATA2[28]), .B2(DATA2[27]), .A(net76578), .ZN(n1302) );
  NOR4_X1 U1293 ( .A1(DATA2[28]), .A2(DATA2[27]), .A3(n1303), .A4(n1185), .ZN(
        n1301) );
  OR2_X1 U1294 ( .A1(DATA2[29]), .A2(DATA2[30]), .ZN(n1185) );
  NOR3_X1 U1295 ( .A1(n1581), .A2(n1580), .A3(n1304), .ZN(n1303) );
  NOR4_X1 U1296 ( .A1(DATA2[26]), .A2(DATA2[25]), .A3(n1305), .A4(n1186), .ZN(
        n1304) );
  AOI22_X1 U1297 ( .A1(net76578), .A2(n1306), .B1(n1670), .B2(n1260), .ZN(
        n1305) );
  OR2_X1 U1298 ( .A1(n1307), .A2(n1308), .ZN(n1260) );
  OAI21_X1 U1299 ( .B1(n1645), .B2(n1692), .A(n1309), .ZN(n1308) );
  AOI22_X1 U1300 ( .A1(n357), .A2(n491), .B1(n356), .B2(n376), .ZN(n1309) );
  NAND2_X1 U1301 ( .A1(n1310), .A2(n1311), .ZN(n376) );
  AOI22_X1 U1302 ( .A1(DATA1[8]), .A2(net76071), .B1(DATA1[7]), .B2(n1527), 
        .ZN(n1311) );
  AOI22_X1 U1303 ( .A1(DATA1[10]), .A2(net76091), .B1(DATA1[9]), .B2(net76107), 
        .ZN(n1310) );
  NOR2_X1 U1304 ( .A1(n1693), .A2(n1442), .ZN(n356) );
  NAND2_X1 U1305 ( .A1(n1312), .A2(n1313), .ZN(n491) );
  AOI22_X1 U1306 ( .A1(DATA1[12]), .A2(net76071), .B1(DATA1[11]), .B2(n1527), 
        .ZN(n1313) );
  AOI22_X1 U1307 ( .A1(DATA1[14]), .A2(net76089), .B1(DATA1[13]), .B2(net76107), .ZN(n1312) );
  NOR2_X1 U1308 ( .A1(net74118), .A2(n1442), .ZN(n357) );
  NOR2_X1 U1309 ( .A1(n1695), .A2(n1442), .ZN(n361) );
  NAND2_X1 U1310 ( .A1(n1314), .A2(n1315), .ZN(n498) );
  AOI22_X1 U1311 ( .A1(n1449), .A2(net76069), .B1(n1448), .B2(n1530), .ZN(
        n1315) );
  AOI22_X1 U1312 ( .A1(DATA1[6]), .A2(net76091), .B1(DATA1[5]), .B2(net76778), 
        .ZN(n1314) );
  NAND2_X1 U1313 ( .A1(n1316), .A2(n1317), .ZN(n1307) );
  AOI22_X1 U1314 ( .A1(n1442), .A2(n905), .B1(n405), .B2(n1318), .ZN(n1317) );
  OAI21_X1 U1315 ( .B1(net81902), .B2(n1657), .A(n1319), .ZN(n1318) );
  AOI21_X1 U1316 ( .B1(n1446), .B2(net76087), .A(n1152), .ZN(n1319) );
  NOR2_X1 U1317 ( .A1(n1660), .A2(n1703), .ZN(n1152) );
  NOR2_X1 U1318 ( .A1(net74115), .A2(n1442), .ZN(n405) );
  OAI21_X1 U1319 ( .B1(n1583), .B2(net74118), .A(n1320), .ZN(n905) );
  NAND2_X1 U1320 ( .A1(n562), .A2(n735), .ZN(n1320) );
  NAND2_X1 U1321 ( .A1(n1321), .A2(n1322), .ZN(n735) );
  AOI22_X1 U1322 ( .A1(DATA1[24]), .A2(net76067), .B1(DATA1[23]), .B2(n1528), 
        .ZN(n1322) );
  AOI22_X1 U1323 ( .A1(DATA1[26]), .A2(net76091), .B1(DATA1[25]), .B2(net76107), .ZN(n1321) );
  NOR2_X1 U1324 ( .A1(n1694), .A2(DATA2[2]), .ZN(n562) );
  NOR2_X1 U1325 ( .A1(n1694), .A2(n1696), .ZN(n563) );
  NAND2_X1 U1326 ( .A1(n1323), .A2(n1324), .ZN(n839) );
  AOI22_X1 U1327 ( .A1(DATA1[28]), .A2(net76067), .B1(DATA1[27]), .B2(n1528), 
        .ZN(n1324) );
  AOI22_X1 U1328 ( .A1(DATA1[30]), .A2(net76091), .B1(net76107), .B2(DATA1[29]), .ZN(n1323) );
  AOI22_X1 U1329 ( .A1(n359), .A2(n374), .B1(n456), .B2(n381), .ZN(n1316) );
  NAND2_X1 U1330 ( .A1(n1325), .A2(n1326), .ZN(n381) );
  AOI22_X1 U1331 ( .A1(DATA1[16]), .A2(net76071), .B1(DATA1[15]), .B2(n1530), 
        .ZN(n1326) );
  AOI22_X1 U1332 ( .A1(DATA1[18]), .A2(net76091), .B1(DATA1[17]), .B2(net76107), .ZN(n1325) );
  NOR2_X1 U1333 ( .A1(net74115), .A2(n1687), .ZN(n456) );
  NOR2_X1 U1334 ( .A1(n1439), .A2(DATA2[2]), .ZN(n576) );
  NAND2_X1 U1335 ( .A1(n1327), .A2(n1328), .ZN(n374) );
  AOI22_X1 U1336 ( .A1(DATA1[20]), .A2(net76067), .B1(DATA1[19]), .B2(n1527), 
        .ZN(n1328) );
  AOI22_X1 U1339 ( .A1(DATA1[22]), .A2(net76089), .B1(DATA1[21]), .B2(net76778), .ZN(n1327) );
  NOR2_X1 U1342 ( .A1(n1695), .A2(n1687), .ZN(n359) );
  NOR2_X1 U1343 ( .A1(n1696), .A2(n1439), .ZN(n465) );
  NAND2_X1 U1344 ( .A1(n1142), .A2(n1671), .ZN(n1306) );
  NOR2_X1 U1345 ( .A1(n1684), .A2(n1181), .ZN(n1142) );
  NAND2_X1 U1346 ( .A1(n1329), .A2(n1330), .ZN(n1181) );
  NOR4_X1 U1347 ( .A1(DATA2[18]), .A2(n1430), .A3(n1428), .A4(n1424), .ZN(
        n1330) );
  NOR3_X1 U1348 ( .A1(n1291), .A2(net82738), .A3(n1290), .ZN(n1329) );
  NAND2_X1 U1349 ( .A1(n1331), .A2(net74147), .ZN(n1290) );
  NOR2_X1 U1350 ( .A1(DATA2[17]), .A2(DATA2[16]), .ZN(n1331) );
  NAND2_X1 U1351 ( .A1(n1332), .A2(n1677), .ZN(n1291) );
  NOR2_X1 U1352 ( .A1(n1417), .A2(n1429), .ZN(n1332) );
  NOR2_X1 U1353 ( .A1(n1333), .A2(n1425), .ZN(n1180) );
  OR2_X1 U1354 ( .A1(n1427), .A2(n1401), .ZN(n1333) );
  NAND2_X1 U1355 ( .A1(net76578), .A2(n1186), .ZN(n1178) );
  NAND2_X1 U1356 ( .A1(n1334), .A2(n1289), .ZN(n1186) );
  NOR2_X1 U1357 ( .A1(n1335), .A2(DATA2[22]), .ZN(n1289) );
  OR2_X1 U1358 ( .A1(DATA2[24]), .A2(DATA2[23]), .ZN(n1335) );
  NOR2_X1 U1359 ( .A1(DATA2[21]), .A2(DATA2[20]), .ZN(n1334) );
  OAI21_X1 U1360 ( .B1(DATA2[26]), .B2(DATA2[25]), .A(net76578), .ZN(n1336) );
  AOI22_X1 U1361 ( .A1(n1274), .A2(n251), .B1(net81160), .B2(n1277), .ZN(n1295) );
  XNOR2_X1 U1362 ( .A(net76759), .B(N1568), .ZN(n1277) );
  AOI21_X1 U1365 ( .B1(net76759), .B2(N1573), .A(n1337), .ZN(n1274) );
  NOR2_X1 U1366 ( .A1(n1538), .A2(net76759), .ZN(n1337) );
  XNOR2_X1 U1371 ( .A(net83443), .B(net94830), .ZN(n320) );
  NOR2_X1 U1372 ( .A1(n1114), .A2(net76566), .ZN(n1208) );
  NAND2_X1 U1374 ( .A1(net83262), .A2(net74079), .ZN(n1191) );
  AOI22_X1 U1153 ( .A1(net82966), .A2(n1204), .B1(net84449), .B2(n306), .ZN(
        n1199) );
  OAI21_X1 U436 ( .B1(n302), .B2(n528), .A(net82966), .ZN(n527) );
  AOI22_X1 U1161 ( .A1(n1145), .A2(net82966), .B1(n315), .B2(n1208), .ZN(n1207) );
  AOI21_X1 U794 ( .B1(n902), .B2(net76161), .A(n1391), .ZN(n901) );
  NAND2_X1 U844 ( .A1(n1393), .A2(net76167), .ZN(n942) );
  NAND2_X1 U818 ( .A1(n1392), .A2(net76167), .ZN(n916) );
  NAND2_X1 U267 ( .A1(n287), .A2(n286), .ZN(n255) );
  NAND2_X1 U1121 ( .A1(n302), .A2(net76759), .ZN(n1166) );
  NOR4_X1 U1242 ( .A1(n1265), .A2(net94964), .A3(net83262), .A4(ALU_OPCODE[4]), 
        .ZN(n1264) );
  OAI33_X1 U1113 ( .A1(n1163), .A2(n1710), .A3(net74084), .B1(n1164), .B2(
        ALU_OPCODE[4]), .B3(net84501), .ZN(n1161) );
  NOR2_X1 U1165 ( .A1(net82584), .A2(net82899), .ZN(n301) );
  AOI21_X1 U254 ( .B1(n249), .B2(n250), .A(net83235), .ZN(n1339) );
  OAI21_X1 U1143 ( .B1(net84454), .B2(net76759), .A(net82953), .ZN(n1190) );
  AOI21_X1 U1142 ( .B1(n1190), .B2(n1191), .A(n1368), .ZN(n1187) );
  OAI21_X1 U1244 ( .B1(n1266), .B2(n1267), .A(net82767), .ZN(n1265) );
  OAI21_X1 U283 ( .B1(n312), .B2(net77211), .A(n313), .ZN(n305) );
  AOI21_X1 U1139 ( .B1(n1187), .B2(n1155), .A(n1188), .ZN(n1160) );
  NAND2_X1 U1124 ( .A1(N2010), .A2(n1174), .ZN(n1173) );
  NAND2_X1 U1112 ( .A1(n1157), .A2(N2010), .ZN(n1162) );
  OAI21_X1 U1111 ( .B1(n1161), .B2(n1160), .A(n1162), .ZN(NEG) );
  NOR3_X1 U1120 ( .A1(net74299), .A2(net83262), .A3(net76573), .ZN(n1168) );
  OAI21_X1 U291 ( .B1(DATA2[31]), .B2(N2010), .A(n323), .ZN(n322) );
  OR2_X1 U1373 ( .A1(n1191), .A2(net77259), .ZN(n1114) );
  OAI21_X1 U1222 ( .B1(net77259), .B2(n1252), .A(n1158), .ZN(n1249) );
  NOR3_X1 U1277 ( .A1(net74077), .A2(net76573), .A3(n1276), .ZN(n1292) );
  OAI21_X1 U1118 ( .B1(net76759), .B2(n1367), .A(net74077), .ZN(n1170) );
  OAI21_X1 U1117 ( .B1(n1168), .B2(n1169), .A(n1170), .ZN(n1167) );
  NOR3_X1 U527 ( .A1(net74128), .A2(net74244), .A3(net74115), .ZN(n651) );
  NOR4_X1 U526 ( .A1(n648), .A2(n649), .A3(n650), .A4(n651), .ZN(n647) );
  AOI22_X1 U540 ( .A1(n512), .A2(n530), .B1(n514), .B2(n513), .ZN(n644) );
  AOI22_X1 U539 ( .A1(net74123), .A2(n666), .B1(net74124), .B2(n524), .ZN(n645) );
  AOI21_X1 U998 ( .B1(n1070), .B2(net76161), .A(n1362), .ZN(n1060) );
  NAND2_X1 U538 ( .A1(N1637), .A2(net76177), .ZN(n665) );
  AOI22_X1 U505 ( .A1(n272), .A2(net76163), .B1(net76554), .B2(n273), .ZN(n619) );
  AOI22_X1 U524 ( .A1(n273), .A2(net76163), .B1(net76555), .B2(n274), .ZN(n643) );
  NOR3_X1 U1110 ( .A1(n528), .A2(n302), .A3(n1159), .ZN(n1153) );
  OAI21_X1 U1106 ( .B1(n1153), .B2(net83235), .A(n526), .ZN(n362) );
  AOI22_X1 U523 ( .A1(N1638), .A2(net76177), .B1(N2007), .B2(net76505), .ZN(
        n620) );
  NAND2_X1 U422 ( .A1(net82056), .A2(net76165), .ZN(n290) );
  NOR2_X1 U1237 ( .A1(net76759), .A2(ALU_OPCODE[5]), .ZN(n252) );
  AOI21_X1 U256 ( .B1(net81160), .B2(n252), .A(n254), .ZN(n249) );
  AOI21_X1 U1241 ( .B1(n1263), .B2(n1725), .A(n1264), .ZN(n1262) );
  AOI22_X1 U432 ( .A1(net76089), .A2(DATA1[28]), .B1(net76781), .B2(DATA1[29]), 
        .ZN(n516) );
  AOI21_X1 U479 ( .B1(DATA1[29]), .B2(net76069), .A(n591), .ZN(n590) );
  AOI21_X1 U968 ( .B1(net76069), .B2(DATA1[30]), .A(n1049), .ZN(n1030) );
  AOI21_X1 U431 ( .B1(DATA1[30]), .B2(net76069), .A(n519), .ZN(n517) );
  NAND2_X1 U430 ( .A1(n516), .A2(n517), .ZN(n515) );
  AOI22_X1 U429 ( .A1(n512), .A2(n513), .B1(n514), .B2(n515), .ZN(n511) );
  OAI21_X1 U428 ( .B1(n510), .B2(net74147), .A(n511), .ZN(n504) );
  OAI21_X1 U1109 ( .B1(n1340), .B2(net83605), .A(n1158), .ZN(n1156) );
  NOR4_X1 U1368 ( .A1(net83262), .A2(net82953), .A3(n1340), .A4(net83235), 
        .ZN(n1338) );
  NOR2_X1 U1367 ( .A1(n1208), .A2(n1338), .ZN(n363) );
  NAND2_X1 U424 ( .A1(net77226), .A2(net76165), .ZN(n501) );
  OAI21_X1 U1126 ( .B1(n904), .B2(n1175), .A(net74295), .ZN(n509) );
  NAND2_X1 U3 ( .A1(net84499), .A2(n1721), .ZN(net77226) );
  NAND2_X1 U10 ( .A1(n1196), .A2(n509), .ZN(net94967) );
  NAND2_X1 U11 ( .A1(N2010), .A2(net83361), .ZN(net82779) );
  NOR2_X1 U12 ( .A1(net83235), .A2(n1714), .ZN(net83361) );
  NOR2_X1 U14 ( .A1(net82884), .A2(n1714), .ZN(net84501) );
  INV_X1 U15 ( .A(n1112), .ZN(n1194) );
  INV_X1 U17 ( .A(net83235), .ZN(net82966) );
  NAND2_X1 U18 ( .A1(net74087), .A2(net82966), .ZN(net94971) );
  NAND2_X1 U20 ( .A1(N1641), .A2(net76177), .ZN(n1238) );
  INV_X2 U21 ( .A(n1198), .ZN(net76177) );
  NAND2_X1 U26 ( .A1(net94971), .A2(n1244), .ZN(n1196) );
  AOI21_X1 U28 ( .B1(n1021), .B2(n1196), .A(n1732), .ZN(n1020) );
  NAND2_X1 U29 ( .A1(n1237), .A2(n1208), .ZN(n1244) );
  NOR2_X1 U30 ( .A1(net94830), .A2(net83422), .ZN(n1237) );
  INV_X1 U31 ( .A(ALU_OPCODE[0]), .ZN(net94830) );
  INV_X1 U33 ( .A(n509), .ZN(net74299) );
  NAND2_X1 U34 ( .A1(n501), .A2(net82927), .ZN(OUTALU[30]) );
  OR2_X1 U35 ( .A1(n1341), .A2(net76169), .ZN(net82927) );
  CLKBUF_X1 U36 ( .A(net74099), .Z(net76169) );
  INV_X1 U37 ( .A(net76553), .ZN(net74099) );
  CLKBUF_X1 U38 ( .A(n363), .Z(net76553) );
  INV_X1 U39 ( .A(n284), .ZN(n1341) );
  CLKBUF_X1 U40 ( .A(net74099), .Z(net76165) );
  CLKBUF_X1 U41 ( .A(n363), .Z(net76554) );
  CLKBUF_X1 U42 ( .A(n363), .Z(net76555) );
  INV_X1 U43 ( .A(n320), .ZN(n1340) );
  INV_X1 U45 ( .A(net74079), .ZN(net82953) );
  INV_X1 U46 ( .A(ALU_OPCODE[2]), .ZN(net74079) );
  INV_X1 U50 ( .A(net84454), .ZN(net83262) );
  CLKBUF_X1 U51 ( .A(net82743), .Z(net84454) );
  NOR2_X1 U52 ( .A1(net84454), .A2(net83605), .ZN(net84449) );
  INV_X1 U53 ( .A(ALU_OPCODE[5]), .ZN(net82743) );
  NOR2_X1 U55 ( .A1(net83605), .A2(net82743), .ZN(n254) );
  NOR3_X1 U56 ( .A1(net77226), .A2(n288), .A3(n1712), .ZN(n287) );
  INV_X1 U63 ( .A(n504), .ZN(net77228) );
  INV_X1 U75 ( .A(n1704), .ZN(net76091) );
  NAND2_X1 U77 ( .A1(net94830), .A2(n1172), .ZN(net83343) );
  INV_X1 U79 ( .A(ALU_OPCODE[1]), .ZN(net74076) );
  NAND2_X1 U80 ( .A1(net77211), .A2(ALU_OPCODE[4]), .ZN(net83422) );
  NOR2_X1 U81 ( .A1(net83422), .A2(net83343), .ZN(net77192) );
  INV_X1 U84 ( .A(ALU_OPCODE[6]), .ZN(net77211) );
  CLKBUF_X1 U85 ( .A(ALU_OPCODE[3]), .Z(net76566) );
  NAND2_X1 U87 ( .A1(ALU_OPCODE[2]), .A2(ALU_OPCODE[1]), .ZN(net83605) );
  CLKBUF_X1 U88 ( .A(ALU_OPCODE[1]), .Z(net83443) );
  OR2_X1 U89 ( .A1(ALU_OPCODE[6]), .A2(ALU_OPCODE[4]), .ZN(net82899) );
  NAND2_X1 U94 ( .A1(n456), .A2(n1347), .ZN(n925) );
  NAND2_X1 U95 ( .A1(n1348), .A2(n290), .ZN(OUTALU[31]) );
  NOR2_X1 U96 ( .A1(net76493), .A2(net76578), .ZN(n1349) );
  AOI21_X1 U99 ( .B1(n1351), .B2(net76578), .A(n1352), .ZN(net145611) );
  NAND2_X1 U106 ( .A1(n1357), .A2(net76159), .ZN(n1351) );
  OAI21_X1 U107 ( .B1(n1349), .B2(net76487), .A(DATA2[31]), .ZN(n1358) );
  NAND2_X1 U109 ( .A1(n534), .A2(n1347), .ZN(net145613) );
  NAND2_X1 U110 ( .A1(net74130), .A2(n535), .ZN(net145612) );
  NAND2_X1 U112 ( .A1(n405), .A2(n402), .ZN(n1359) );
  NAND2_X1 U114 ( .A1(net145680), .A2(net76555), .ZN(n1348) );
  NAND2_X1 U116 ( .A1(n620), .A2(n1737), .ZN(n272) );
  CLKBUF_X1 U117 ( .A(n362), .Z(net76505) );
  AOI22_X1 U119 ( .A1(N1638), .A2(net76177), .B1(N2007), .B2(net76505), .ZN(
        net107648) );
  CLKBUF_X1 U120 ( .A(n362), .Z(net76506) );
  CLKBUF_X1 U121 ( .A(n362), .Z(net76507) );
  NOR2_X1 U123 ( .A1(net84454), .A2(net74079), .ZN(n302) );
  NOR3_X1 U125 ( .A1(n1361), .A2(n273), .A3(n271), .ZN(n270) );
  OR2_X1 U127 ( .A1(n272), .A2(n274), .ZN(n1361) );
  INV_X1 U129 ( .A(net82738), .ZN(n1362) );
  CLKBUF_X1 U130 ( .A(DATA2[11]), .Z(net82738) );
  NAND2_X1 U131 ( .A1(n1723), .A2(n1706), .ZN(n1365) );
  INV_X1 U134 ( .A(n522), .ZN(net74124) );
  INV_X1 U135 ( .A(n747), .ZN(net74123) );
  INV_X1 U138 ( .A(n576), .ZN(net74115) );
  INV_X1 U140 ( .A(n926), .ZN(net74244) );
  NAND2_X1 U141 ( .A1(n1167), .A2(net83745), .ZN(n1164) );
  INV_X1 U142 ( .A(n314), .ZN(net74077) );
  NAND2_X1 U144 ( .A1(net82953), .A2(net77259), .ZN(n1367) );
  CLKBUF_X1 U147 ( .A(net74076), .Z(net77259) );
  CLKBUF_X1 U149 ( .A(net94830), .Z(net76759) );
  INV_X1 U153 ( .A(N2010), .ZN(net82884) );
  OR2_X1 U156 ( .A1(net82884), .A2(n1166), .ZN(net83745) );
  NAND2_X1 U157 ( .A1(net83235), .A2(n1369), .ZN(n1188) );
  NAND2_X1 U158 ( .A1(n1208), .A2(n1736), .ZN(n1369) );
  CLKBUF_X1 U161 ( .A(ALU_OPCODE[6]), .Z(net82767) );
  INV_X1 U162 ( .A(n1192), .ZN(n1368) );
  NAND2_X1 U165 ( .A1(net94830), .A2(n251), .ZN(n250) );
  OR2_X1 U166 ( .A1(net82899), .A2(net76566), .ZN(net83235) );
  CLKBUF_X1 U167 ( .A(net82899), .Z(net84429) );
  INV_X1 U168 ( .A(ALU_OPCODE[4]), .ZN(net74084) );
  NOR2_X1 U169 ( .A1(n284), .A2(n1371), .ZN(n1406) );
  NAND2_X1 U170 ( .A1(n1419), .A2(n278), .ZN(n1371) );
  NAND2_X1 U172 ( .A1(net95157), .A2(n1711), .ZN(n1404) );
  INV_X1 U176 ( .A(n741), .ZN(n1379) );
  INV_X1 U180 ( .A(n1375), .ZN(n714) );
  OR2_X1 U187 ( .A1(n1383), .A2(n686), .ZN(n274) );
  NAND2_X1 U188 ( .A1(n1724), .A2(n1705), .ZN(n1383) );
  INV_X1 U190 ( .A(n696), .ZN(n1390) );
  INV_X1 U205 ( .A(n894), .ZN(n1392) );
  INV_X1 U206 ( .A(n915), .ZN(n1393) );
  NAND2_X1 U207 ( .A1(net84505), .A2(n1399), .ZN(n288) );
  OR2_X1 U208 ( .A1(net84507), .A2(n1398), .ZN(n1399) );
  NAND2_X1 U211 ( .A1(net82651), .A2(n1733), .ZN(net82056) );
  OR2_X1 U213 ( .A1(n1391), .A2(n510), .ZN(n1395) );
  INV_X1 U214 ( .A(DATA2[16]), .ZN(n1391) );
  INV_X1 U216 ( .A(n405), .ZN(net74119) );
  CLKBUF_X1 U220 ( .A(DATA2[6]), .Z(n1401) );
  NAND2_X1 U223 ( .A1(n1715), .A2(n596), .ZN(n271) );
  INV_X1 U225 ( .A(net81160), .ZN(net94951) );
  NOR2_X1 U226 ( .A1(net76573), .A2(net94906), .ZN(n1144) );
  NOR2_X1 U228 ( .A1(net81160), .A2(n314), .ZN(n1253) );
  OAI21_X1 U231 ( .B1(net74079), .B2(ALU_OPCODE[0]), .A(net94951), .ZN(
        net94964) );
  CLKBUF_X1 U236 ( .A(DATA2[8]), .Z(n1429) );
  CLKBUF_X1 U237 ( .A(ALU_OPCODE[0]), .Z(net76573) );
  CLKBUF_X1 U238 ( .A(DATA1[0]), .Z(n1444) );
  NAND2_X1 U245 ( .A1(N2011), .A2(n1408), .ZN(net84505) );
  INV_X1 U246 ( .A(net82941), .ZN(net84507) );
  NAND2_X1 U248 ( .A1(N2010), .A2(n1418), .ZN(net84496) );
  NOR2_X1 U249 ( .A1(n1717), .A2(n1414), .ZN(net84497) );
  CLKBUF_X1 U255 ( .A(DATA2[4]), .Z(n1442) );
  CLKBUF_X1 U288 ( .A(DATA1[1]), .Z(n1411) );
  OR2_X1 U423 ( .A1(n322), .A2(net77259), .ZN(n319) );
  OR2_X1 U426 ( .A1(n321), .A2(net74092), .ZN(n1413) );
  NAND2_X1 U427 ( .A1(n1413), .A2(net74309), .ZN(n317) );
  NOR2_X1 U437 ( .A1(n747), .A2(net83387), .ZN(n1414) );
  INV_X1 U439 ( .A(n524), .ZN(net83387) );
  OR2_X1 U441 ( .A1(net82652), .A2(n1431), .ZN(n1415) );
  NAND2_X1 U442 ( .A1(N2011), .A2(n1415), .ZN(net82651) );
  INV_X1 U466 ( .A(n1199), .ZN(net82652) );
  INV_X1 U486 ( .A(n1200), .ZN(n1431) );
  INV_X1 U536 ( .A(n1698), .ZN(n1416) );
  CLKBUF_X1 U546 ( .A(DATA2[9]), .Z(n1417) );
  OR2_X1 U568 ( .A1(net82924), .A2(net82925), .ZN(n1418) );
  NOR3_X1 U746 ( .A1(n283), .A2(n282), .A3(n1553), .ZN(n1419) );
  CLKBUF_X1 U932 ( .A(DATA2[1]), .Z(n1420) );
  OR2_X1 U1119 ( .A1(net83262), .A2(net82953), .ZN(n1421) );
  NAND2_X1 U1140 ( .A1(n316), .A2(n1421), .ZN(n294) );
  OR2_X1 U1146 ( .A1(net82942), .A2(net76165), .ZN(net82941) );
  INV_X1 U1147 ( .A(net82933), .ZN(net82942) );
  OR2_X1 U1154 ( .A1(n289), .A2(net76169), .ZN(net82933) );
  INV_X1 U1155 ( .A(n526), .ZN(net82924) );
  INV_X1 U1163 ( .A(n527), .ZN(net82925) );
  NAND2_X1 U1209 ( .A1(n1716), .A2(n569), .ZN(n284) );
  INV_X1 U1214 ( .A(net84429), .ZN(n306) );
  CLKBUF_X1 U1215 ( .A(DATA2[12]), .Z(n1424) );
  CLKBUF_X1 U1225 ( .A(DATA2[5]), .Z(n1425) );
  CLKBUF_X1 U1243 ( .A(DATA2[10]), .Z(n1426) );
  CLKBUF_X1 U1251 ( .A(DATA2[13]), .Z(n1428) );
  CLKBUF_X1 U1279 ( .A(DATA2[14]), .Z(n1430) );
  OR2_X1 U1337 ( .A1(net94830), .A2(net83262), .ZN(net82724) );
  CLKBUF_X1 U1363 ( .A(n352), .Z(n1434) );
  INV_X1 U1364 ( .A(n1195), .ZN(net82057) );
  INV_X1 U1369 ( .A(net76566), .ZN(net82584) );
  NOR2_X1 U1370 ( .A1(n1404), .A2(n255), .ZN(ZERO) );
  INV_X1 U1375 ( .A(net76501), .ZN(net74121) );
  INV_X1 U1378 ( .A(n658), .ZN(n1685) );
  INV_X1 U1379 ( .A(n411), .ZN(n1662) );
  CLKBUF_X1 U1380 ( .A(n514), .Z(net76501) );
  CLKBUF_X1 U1381 ( .A(net76149), .Z(net76147) );
  CLKBUF_X1 U1382 ( .A(n512), .Z(net76479) );
  INV_X1 U1383 ( .A(n397), .ZN(n1689) );
  INV_X1 U1386 ( .A(n661), .ZN(n1664) );
  CLKBUF_X1 U1387 ( .A(net76778), .Z(net76781) );
  CLKBUF_X1 U1388 ( .A(net76107), .Z(net76778) );
  INV_X1 U1389 ( .A(n534), .ZN(net74120) );
  INV_X1 U1390 ( .A(n628), .ZN(n1688) );
  INV_X1 U1392 ( .A(n819), .ZN(n1567) );
  INV_X1 U1393 ( .A(n359), .ZN(net74135) );
  INV_X1 U1394 ( .A(n614), .ZN(n1647) );
  INV_X1 U1395 ( .A(n436), .ZN(n1565) );
  INV_X1 U1397 ( .A(n1704), .ZN(net76089) );
  INV_X1 U1399 ( .A(n1704), .ZN(net76087) );
  INV_X1 U1401 ( .A(net81902), .ZN(net76107) );
  INV_X1 U1402 ( .A(n1509), .ZN(n1695) );
  INV_X1 U1403 ( .A(n456), .ZN(net74133) );
  INV_X1 U1404 ( .A(n964), .ZN(n1682) );
  INV_X1 U1405 ( .A(n415), .ZN(n1681) );
  INV_X1 U1406 ( .A(n361), .ZN(n1692) );
  INV_X1 U1407 ( .A(n333), .ZN(n1679) );
  INV_X1 U1408 ( .A(n492), .ZN(n1680) );
  INV_X1 U1409 ( .A(n344), .ZN(n1571) );
  INV_X1 U1410 ( .A(n445), .ZN(n1683) );
  INV_X1 U1411 ( .A(n519), .ZN(net74307) );
  INV_X1 U1412 ( .A(n781), .ZN(n1654) );
  INV_X1 U1413 ( .A(n578), .ZN(n1566) );
  INV_X1 U1414 ( .A(n723), .ZN(n1659) );
  INV_X1 U1415 ( .A(n462), .ZN(n1656) );
  INV_X1 U1424 ( .A(net76535), .ZN(net74118) );
  INV_X1 U1425 ( .A(n650), .ZN(net74292) );
  INV_X1 U1427 ( .A(n388), .ZN(n1686) );
  INV_X1 U1428 ( .A(n601), .ZN(n1544) );
  INV_X1 U1429 ( .A(n684), .ZN(n1562) );
  INV_X1 U1430 ( .A(n1520), .ZN(n1691) );
  INV_X1 U1431 ( .A(n407), .ZN(n1575) );
  INV_X1 U1432 ( .A(n419), .ZN(n1570) );
  INV_X1 U1433 ( .A(n941), .ZN(n1559) );
  INV_X1 U1434 ( .A(n324), .ZN(n1554) );
  INV_X1 U1435 ( .A(n966), .ZN(n1539) );
  INV_X1 U1436 ( .A(n736), .ZN(n1548) );
  INV_X1 U1437 ( .A(N1576), .ZN(n1535) );
  INV_X1 U1438 ( .A(n1029), .ZN(n1563) );
  INV_X1 U1439 ( .A(n1434), .ZN(n1690) );
  INV_X1 U1440 ( .A(n1703), .ZN(net76069) );
  INV_X1 U1441 ( .A(n1703), .ZN(net76071) );
  INV_X1 U1442 ( .A(n1703), .ZN(net76067) );
  INV_X1 U1443 ( .A(n546), .ZN(n1665) );
  INV_X1 U1444 ( .A(n1435), .ZN(n1527) );
  INV_X1 U1445 ( .A(n1435), .ZN(n1528) );
  INV_X1 U1447 ( .A(n1435), .ZN(n1530) );
  INV_X1 U1448 ( .A(n370), .ZN(n1560) );
  INV_X1 U1449 ( .A(n428), .ZN(n1644) );
  INV_X1 U1450 ( .A(n735), .ZN(n1589) );
  INV_X1 U1451 ( .A(net76505), .ZN(net74162) );
  INV_X1 U1452 ( .A(n283), .ZN(n1552) );
  INV_X1 U1453 ( .A(n1511), .ZN(n1693) );
  INV_X1 U1454 ( .A(n1176), .ZN(net74295) );
  INV_X1 U1455 ( .A(n350), .ZN(n1701) );
  INV_X1 U1456 ( .A(n703), .ZN(net74128) );
  INV_X1 U1457 ( .A(n582), .ZN(n1700) );
  CLKBUF_X1 U1458 ( .A(net76061), .Z(net76063) );
  INV_X1 U1459 ( .A(n905), .ZN(n1582) );
  INV_X1 U1460 ( .A(n472), .ZN(n1612) );
  INV_X1 U1462 ( .A(n387), .ZN(n1564) );
  INV_X1 U1463 ( .A(n636), .ZN(n1630) );
  INV_X1 U1464 ( .A(n486), .ZN(n1569) );
  INV_X1 U1465 ( .A(n547), .ZN(n1577) );
  INV_X1 U1466 ( .A(n808), .ZN(n1568) );
  INV_X1 U1467 ( .A(n610), .ZN(n1618) );
  CLKBUF_X1 U1468 ( .A(net76061), .Z(net76065) );
  INV_X1 U1469 ( .A(n418), .ZN(n1555) );
  INV_X1 U1470 ( .A(n381), .ZN(n1615) );
  INV_X1 U1471 ( .A(n713), .ZN(net74130) );
  CLKBUF_X1 U1474 ( .A(n465), .Z(n1509) );
  CLKBUF_X1 U1481 ( .A(n357), .Z(n1517) );
  INV_X1 U1482 ( .A(n408), .ZN(n1619) );
  INV_X1 U1483 ( .A(n360), .ZN(n1576) );
  INV_X1 U1484 ( .A(n336), .ZN(n1597) );
  INV_X1 U1485 ( .A(n285), .ZN(n1553) );
  INV_X1 U1486 ( .A(n774), .ZN(n1585) );
  INV_X1 U1487 ( .A(n1068), .ZN(n1578) );
  INV_X1 U1488 ( .A(n800), .ZN(n1648) );
  INV_X1 U1489 ( .A(n473), .ZN(n1633) );
  CLKBUF_X1 U1490 ( .A(n356), .Z(n1520) );
  INV_X1 U1491 ( .A(n1145), .ZN(net74089) );
  INV_X1 U1494 ( .A(n438), .ZN(n1609) );
  INV_X1 U1495 ( .A(n409), .ZN(n1605) );
  INV_X1 U1496 ( .A(n460), .ZN(n1587) );
  INV_X1 U1497 ( .A(n437), .ZN(n1622) );
  INV_X1 U1498 ( .A(n498), .ZN(n1645) );
  INV_X1 U1499 ( .A(n839), .ZN(n1583) );
  INV_X1 U1500 ( .A(n659), .ZN(n1632) );
  INV_X1 U1501 ( .A(n639), .ZN(n1640) );
  INV_X1 U1502 ( .A(n635), .ZN(n1623) );
  INV_X1 U1503 ( .A(n491), .ZN(n1626) );
  INV_X1 U1504 ( .A(n682), .ZN(n1634) );
  INV_X1 U1505 ( .A(n346), .ZN(n1637) );
  INV_X1 U1506 ( .A(n374), .ZN(n1602) );
  CLKBUF_X1 U1507 ( .A(n563), .Z(net76535) );
  INV_X1 U1508 ( .A(n1027), .ZN(n1663) );
  INV_X1 U1509 ( .A(n611), .ZN(n1628) );
  INV_X1 U1510 ( .A(n1182), .ZN(n1579) );
  INV_X1 U1511 ( .A(n751), .ZN(n1584) );
  INV_X1 U1512 ( .A(n733), .ZN(n1594) );
  INV_X1 U1513 ( .A(N1979), .ZN(n1658) );
  INV_X1 U1514 ( .A(n435), .ZN(n1639) );
  INV_X1 U1515 ( .A(n332), .ZN(n1598) );
  INV_X1 U1516 ( .A(n1126), .ZN(n1596) );
  INV_X1 U1517 ( .A(n1063), .ZN(n1557) );
  INV_X1 U1518 ( .A(n510), .ZN(net74095) );
  CLKBUF_X1 U1519 ( .A(net74099), .Z(net76163) );
  CLKBUF_X1 U1520 ( .A(net74099), .Z(net76167) );
  CLKBUF_X1 U1521 ( .A(net76487), .Z(net76488) );
  INV_X1 U1522 ( .A(n271), .ZN(net74296) );
  INV_X1 U1523 ( .A(n530), .ZN(net74227) );
  INV_X1 U1524 ( .A(n292), .ZN(n1556) );
  INV_X1 U1525 ( .A(n281), .ZN(n1543) );
  INV_X1 U1526 ( .A(n276), .ZN(n1549) );
  INV_X1 U1527 ( .A(n998), .ZN(n1558) );
  INV_X1 U1528 ( .A(n983), .ZN(n1572) );
  INV_X1 U1529 ( .A(n264), .ZN(n1547) );
  INV_X1 U1530 ( .A(n1236), .ZN(net74087) );
  INV_X1 U1531 ( .A(N1999), .ZN(n1606) );
  INV_X1 U1532 ( .A(N1998), .ZN(n1610) );
  INV_X1 U1533 ( .A(N1995), .ZN(n1620) );
  INV_X1 U1534 ( .A(n827), .ZN(n1607) );
  INV_X1 U1535 ( .A(N1577), .ZN(n1536) );
  INV_X1 U1536 ( .A(n619), .ZN(net74300) );
  INV_X1 U1537 ( .A(n643), .ZN(net74287) );
  INV_X1 U1538 ( .A(n876), .ZN(OUTALU[16]) );
  INV_X1 U1539 ( .A(n822), .ZN(OUTALU[19]) );
  INV_X1 U1540 ( .A(n858), .ZN(OUTALU[17]) );
  INV_X1 U1541 ( .A(n840), .ZN(OUTALU[18]) );
  INV_X1 U1542 ( .A(N1572), .ZN(n1538) );
  INV_X1 U1543 ( .A(n1251), .ZN(n1537) );
  INV_X1 U1544 ( .A(n1442), .ZN(n1687) );
  INV_X1 U1545 ( .A(n801), .ZN(OUTALU[1]) );
  INV_X1 U1546 ( .A(n724), .ZN(n1641) );
  INV_X1 U1547 ( .A(n1181), .ZN(n1673) );
  INV_X1 U1548 ( .A(n280), .ZN(n1561) );
  INV_X1 U1549 ( .A(n301), .ZN(net74096) );
  INV_X1 U1550 ( .A(DATA1[9]), .ZN(n1636) );
  INV_X1 U1551 ( .A(DATA1[17]), .ZN(n1617) );
  INV_X1 U1552 ( .A(n496), .ZN(n1541) );
  INV_X1 U1553 ( .A(DATA1[11]), .ZN(n1631) );
  INV_X1 U1554 ( .A(DATA1[16]), .ZN(n1621) );
  INV_X1 U1555 ( .A(DATA1[27]), .ZN(n1586) );
  INV_X1 U1556 ( .A(DATA1[26]), .ZN(n1588) );
  INV_X1 U1557 ( .A(DATA1[7]), .ZN(n1642) );
  INV_X1 U1558 ( .A(DATA1[6]), .ZN(n1643) );
  INV_X1 U1559 ( .A(DATA1[28]), .ZN(net74243) );
  INV_X1 U1560 ( .A(DATA1[10]), .ZN(net74191) );
  CLKBUF_X1 U1561 ( .A(n576), .Z(net76542) );
  INV_X1 U1563 ( .A(n376), .ZN(n1635) );
  INV_X1 U1564 ( .A(n485), .ZN(n1649) );
  INV_X1 U1569 ( .A(net77196), .ZN(net74147) );
  INV_X1 U1570 ( .A(n1179), .ZN(n1667) );
  INV_X1 U1571 ( .A(n1444), .ZN(n1660) );
  INV_X1 U1573 ( .A(n1439), .ZN(n1694) );
  CLKBUF_X1 U1574 ( .A(n562), .Z(n1511) );
  INV_X1 U1576 ( .A(n1449), .ZN(n1651) );
  INV_X1 U1577 ( .A(n1448), .ZN(n1652) );
  INV_X1 U1579 ( .A(n1446), .ZN(n1655) );
  INV_X1 U1580 ( .A(n566), .ZN(n1653) );
  INV_X1 U1581 ( .A(DATA1[30]), .ZN(net74249) );
  INV_X1 U1582 ( .A(n1180), .ZN(n1684) );
  INV_X1 U1583 ( .A(DATA1[12]), .ZN(n1629) );
  INV_X1 U1584 ( .A(DATA2[0]), .ZN(n1698) );
  INV_X1 U1585 ( .A(n725), .ZN(n1650) );
  INV_X1 U1586 ( .A(DATA1[22]), .ZN(n1601) );
  INV_X1 U1587 ( .A(n261), .ZN(n1551) );
  INV_X1 U1588 ( .A(DATA1[13]), .ZN(n1627) );
  INV_X1 U1589 ( .A(DATA1[29]), .ZN(net74246) );
  INV_X1 U1590 ( .A(DATA1[5]), .ZN(n1646) );
  INV_X1 U1591 ( .A(DATA1[23]), .ZN(n1599) );
  INV_X1 U1592 ( .A(n1289), .ZN(n1669) );
  OR2_X1 U1593 ( .A1(n1697), .A2(n1416), .ZN(net81902) );
  INV_X1 U1594 ( .A(DATA1[18]), .ZN(n1614) );
  INV_X1 U1595 ( .A(DATA1[14]), .ZN(n1625) );
  INV_X1 U1596 ( .A(DATA1[15]), .ZN(n1624) );
  INV_X1 U1597 ( .A(DATA1[24]), .ZN(n1593) );
  INV_X1 U1598 ( .A(DATA1[19]), .ZN(n1611) );
  INV_X1 U1599 ( .A(n322), .ZN(net74309) );
  INV_X1 U1601 ( .A(N2003), .ZN(n1592) );
  INV_X1 U1602 ( .A(N1997), .ZN(n1613) );
  INV_X1 U1603 ( .A(N1996), .ZN(n1616) );
  INV_X1 U1604 ( .A(N2000), .ZN(n1603) );
  INV_X1 U1605 ( .A(N2004), .ZN(n1590) );
  INV_X1 U1606 ( .A(N2002), .ZN(n1595) );
  INV_X1 U1607 ( .A(N2001), .ZN(n1600) );
  CLKBUF_X1 U1631 ( .A(DATA1[4]), .Z(n1449) );
  INV_X1 U1632 ( .A(n1306), .ZN(n1670) );
  INV_X1 U1633 ( .A(n1154), .ZN(n1699) );
  INV_X1 U1634 ( .A(n829), .ZN(n1608) );
  INV_X1 U1635 ( .A(n1178), .ZN(n1580) );
  INV_X1 U1636 ( .A(DATA1[25]), .ZN(n1591) );
  INV_X1 U1637 ( .A(DATA1[21]), .ZN(n1604) );
  INV_X1 U1638 ( .A(DATA1[8]), .ZN(n1638) );
  INV_X1 U1639 ( .A(n425), .ZN(n1573) );
  OR2_X1 U1640 ( .A1(n1420), .A2(n1416), .ZN(n1435) );
  INV_X1 U1641 ( .A(n393), .ZN(n1574) );
  INV_X1 U1652 ( .A(n1411), .ZN(n1657) );
  INV_X1 U1654 ( .A(n1420), .ZN(n1697) );
  INV_X1 U1655 ( .A(DATA2[2]), .ZN(n1696) );
  INV_X1 U1656 ( .A(n310), .ZN(n1702) );
  INV_X1 U1669 ( .A(DATA2[19]), .ZN(n1671) );
  CLKBUF_X1 U1676 ( .A(DATA1[2]), .Z(n1446) );
  CLKBUF_X1 U1677 ( .A(DATA2[3]), .Z(n1439) );
  INV_X1 U1682 ( .A(n1426), .ZN(n1677) );
  INV_X1 U1683 ( .A(n1336), .ZN(n1581) );
  INV_X1 U1684 ( .A(n1275), .ZN(n1661) );
  INV_X1 U1687 ( .A(n1424), .ZN(n1676) );
  INV_X1 U1688 ( .A(n1430), .ZN(n1675) );
  INV_X1 U1689 ( .A(DATA2[18]), .ZN(n1672) );
  INV_X1 U1690 ( .A(DATA2[24]), .ZN(n1668) );
  INV_X1 U1691 ( .A(n1417), .ZN(n1678) );
  INV_X1 U1692 ( .A(DATA2[17]), .ZN(n1674) );
  INV_X1 U1693 ( .A(n302), .ZN(net74092) );
  CLKBUF_X1 U1695 ( .A(DATA2[15]), .Z(net77196) );
  CLKBUF_X1 U1696 ( .A(net74099), .Z(net76171) );
  CLKBUF_X1 U1697 ( .A(net76159), .Z(net76161) );
  ALU_N32_DW01_cmp6_0 r167 ( .A({net76578, DATA1[30:5], n1449, n1448, n1446, 
        n1411, n1444}), .B({DATA2[31:16], net77196, n1430, n1428, n1424, 
        net82738, n1426, n1417, n1429, n1427, n1401, n1425, n1442, n1439, 
        DATA2[2], n1420, DATA2[0]}), .TC(1'b1), .LE(N1572), .GE(N1573) );
  ALU_N32_DW01_cmp6_1 r166 ( .A({net76578, DATA1[30:5], n1449, n1448, n1446, 
        n1411, n1444}), .B({DATA2[31:16], net77196, n1430, n1428, n1424, 
        net82738, n1426, n1417, n1429, n1427, n1401, n1425, n1442, n1439, 
        DATA2[2], n1420, n1416}), .TC(1'b0), .EQ(N1568), .LE(N1576), .GE(N1577) );
  ALU_N32_DW02_mult_0 r79 ( .A(DATA1[15:0]), .B(DATA2[15:0]), .TC(\U2/U1/Z_0 ), 
        .PRODUCT({N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, 
        N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, 
        N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, 
        N1613, N1612, N1611, N1610}) );
  ALU_N32_DW01_addsub_2 r170 ( .A({1'b0, net76578, DATA1[30:5], n1449, n1448, 
        n1446, n1411, n1444}), .B({1'b0, DATA2[31:16], net77196, n1430, n1428, 
        n1424, net82738, n1426, n1417, n1429, n1427, n1401, n1425, n1442, 
        n1439, DATA2[2:0]}), .CI(1'b0), .ADD_SUB(n1339), .SUM({N2011, N2010, 
        N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, 
        N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, 
        N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, 
        N1979}) );
  OR2_X1 U2 ( .A1(n1698), .A2(n1420), .ZN(n1703) );
  OR2_X1 U4 ( .A1(n1697), .A2(n1698), .ZN(n1704) );
  AND3_X1 U6 ( .A1(n673), .A2(n670), .A3(n671), .ZN(n1705) );
  AND3_X1 U13 ( .A1(n647), .A2(n644), .A3(n645), .ZN(n1706) );
  AND2_X1 U16 ( .A1(n743), .A2(n744), .ZN(n1707) );
  AND2_X1 U19 ( .A1(n698), .A2(n699), .ZN(n1708) );
  AND2_X1 U22 ( .A1(n259), .A2(n260), .ZN(n1709) );
  AND3_X1 U23 ( .A1(N1641), .A2(n1725), .A3(n321), .ZN(n1710) );
  AND2_X1 U24 ( .A1(n1406), .A2(n1709), .ZN(n1711) );
  OR2_X1 U25 ( .A1(n1393), .A2(n1392), .ZN(n1712) );
  OR4_X1 U27 ( .A1(DATA2[19]), .A2(n1667), .A3(n1185), .A4(n1186), .ZN(n1713)
         );
  OR2_X1 U32 ( .A1(n311), .A2(n1194), .ZN(n1714) );
  AND3_X1 U44 ( .A1(n599), .A2(n597), .A3(n598), .ZN(n1715) );
  AND3_X1 U47 ( .A1(n572), .A2(n570), .A3(n571), .ZN(n1716) );
  NOR2_X1 U48 ( .A1(net74227), .A2(n522), .ZN(n1717) );
  OR3_X1 U49 ( .A1(net74307), .A2(n1207), .A3(net74119), .ZN(n1718) );
  AND2_X1 U54 ( .A1(n756), .A2(n757), .ZN(n1719) );
  AND2_X1 U57 ( .A1(n1730), .A2(net84497), .ZN(n1720) );
  AND2_X1 U58 ( .A1(net84496), .A2(n1720), .ZN(n1721) );
  AND2_X1 U59 ( .A1(n709), .A2(n710), .ZN(n1722) );
  NAND2_X1 U60 ( .A1(N2006), .A2(net76505), .ZN(n1723) );
  NAND2_X1 U61 ( .A1(N2005), .A2(net76507), .ZN(n1724) );
  CLKBUF_X1 U62 ( .A(n1172), .Z(n1725) );
  OR2_X1 U64 ( .A1(net74162), .A2(n1592), .ZN(n1726) );
  NAND2_X1 U65 ( .A1(n731), .A2(n1726), .ZN(n730) );
  AND2_X1 U66 ( .A1(ALU_OPCODE[3]), .A2(net82743), .ZN(n1172) );
  OR2_X1 U67 ( .A1(n510), .A2(n1362), .ZN(n1727) );
  NAND2_X1 U68 ( .A1(n1727), .A2(n665), .ZN(n664) );
  OR2_X2 U69 ( .A1(n1365), .A2(n664), .ZN(n273) );
  AND3_X1 U70 ( .A1(n1722), .A2(n1388), .A3(n1708), .ZN(n1728) );
  AND2_X1 U71 ( .A1(n1390), .A2(n1728), .ZN(n276) );
  AND2_X1 U72 ( .A1(n1238), .A2(net112136), .ZN(net84499) );
  OAI21_X2 U73 ( .B1(net83235), .B2(n1108), .A(n1109), .ZN(net76061) );
  CLKBUF_X1 U74 ( .A(DATA1[3]), .Z(n1448) );
  AND2_X1 U76 ( .A1(net74076), .A2(ALU_OPCODE[2]), .ZN(net81160) );
  AND2_X1 U78 ( .A1(net82779), .A2(net94967), .ZN(net112136) );
  CLKBUF_X1 U82 ( .A(DATA2[7]), .Z(n1427) );
  AND2_X1 U83 ( .A1(n1733), .A2(net82933), .ZN(n1398) );
  NAND4_X1 U86 ( .A1(n1719), .A2(n1377), .A3(n1707), .A4(n1379), .ZN(n1375) );
  INV_X1 U90 ( .A(n739), .ZN(n1377) );
  AND2_X1 U91 ( .A1(ALU_OPCODE[2]), .A2(net83443), .ZN(n251) );
  AND2_X1 U92 ( .A1(net77192), .A2(net81160), .ZN(\U2/U1/Z_0 ) );
  NAND4_X1 U93 ( .A1(n1285), .A2(n1286), .A3(n1287), .A4(n1288), .ZN(n1073) );
  AND2_X1 U97 ( .A1(net76542), .A2(n776), .ZN(n775) );
  INV_X1 U98 ( .A(n1358), .ZN(n1352) );
  MUX2_X1 U100 ( .A(net76493), .B(n1353), .S(DATA2[31]), .Z(n1357) );
  INV_X1 U101 ( .A(net76061), .ZN(n1353) );
  INV_X1 U102 ( .A(n1208), .ZN(net94906) );
  AND2_X1 U103 ( .A1(n1359), .A2(n1729), .ZN(n1088) );
  OR2_X1 U104 ( .A1(n652), .A2(net74135), .ZN(n1729) );
  INV_X1 U105 ( .A(n652), .ZN(n1347) );
  INV_X1 U108 ( .A(n1196), .ZN(net74101) );
  INV_X1 U111 ( .A(net76578), .ZN(net74263) );
  AND2_X1 U113 ( .A1(n588), .A2(n361), .ZN(n587) );
  AND2_X1 U115 ( .A1(n592), .A2(n1520), .ZN(n585) );
  INV_X1 U118 ( .A(net76487), .ZN(net76159) );
  INV_X1 U122 ( .A(net76493), .ZN(net76149) );
  AND4_X1 U124 ( .A1(net145611), .A2(net145612), .A3(net145613), .A4(net77228), 
        .ZN(n1730) );
  INV_X1 U126 ( .A(net94964), .ZN(n1206) );
  AND2_X1 U128 ( .A1(n1415), .A2(net82941), .ZN(n1408) );
  OR2_X1 U132 ( .A1(n1731), .A2(n850), .ZN(n1354) );
  AND2_X1 U133 ( .A1(n563), .A2(n1347), .ZN(n1731) );
  AND2_X1 U136 ( .A1(DATA1[10]), .A2(n1022), .ZN(n1732) );
  INV_X1 U137 ( .A(n1354), .ZN(n564) );
  NAND3_X1 U139 ( .A1(net84499), .A2(net84530), .A3(n1730), .ZN(net145680) );
  AND2_X1 U143 ( .A1(net84496), .A2(net84497), .ZN(net84530) );
  AND3_X1 U145 ( .A1(net82057), .A2(n1718), .A3(n1395), .ZN(n1733) );
  AND2_X1 U146 ( .A1(N2010), .A2(n252), .ZN(n1169) );
  NOR2_X1 U148 ( .A1(n1734), .A2(n1735), .ZN(n1157) );
  OR3_X1 U150 ( .A1(net77211), .A2(net82953), .A3(n321), .ZN(n1734) );
  OR3_X1 U151 ( .A1(net76566), .A2(net83262), .A3(ALU_OPCODE[4]), .ZN(n1735)
         );
  AND2_X1 U152 ( .A1(net76573), .A2(net77211), .ZN(n1736) );
  INV_X1 U154 ( .A(net83422), .ZN(n315) );
  NAND4_X1 U155 ( .A1(n802), .A2(n803), .A3(n804), .A4(n805), .ZN(n261) );
  NAND4_X1 U159 ( .A1(n539), .A2(n540), .A3(n541), .A4(n542), .ZN(n283) );
  NAND4_X1 U160 ( .A1(n478), .A2(n479), .A3(n480), .A4(n481), .ZN(n282) );
  NAND4_X1 U163 ( .A1(n422), .A2(n423), .A3(n424), .A4(n1573), .ZN(n280) );
  NAND4_X1 U164 ( .A1(n390), .A2(n391), .A3(n392), .A4(n1574), .ZN(n279) );
  NAND4_X1 U171 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n291) );
  INV_X1 U173 ( .A(n694), .ZN(n1388) );
  AND3_X1 U174 ( .A1(n623), .A2(n621), .A3(n622), .ZN(n1737) );
  NAND3_X1 U175 ( .A1(n1725), .A2(n315), .A3(net81160), .ZN(n1198) );
  AND2_X1 U177 ( .A1(n270), .A2(n269), .ZN(net95157) );
  AND2_X1 U178 ( .A1(n1737), .A2(net107648), .ZN(n1374) );
endmodule


module gen_reg_N32_4 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n103, n110, n111, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n173), .B2(n111), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n110), .A2(data_in[23]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n174), .B2(ld), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[24]), .A2(n111), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n175), .B2(ld), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[25]), .A2(n111), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n176), .B2(ld), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[26]), .A2(n110), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n177), .B2(n111), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[27]), .A2(n110), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n178), .B2(ld), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[28]), .A2(n111), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n110), .A(n143), .ZN(n32) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n111), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n111), .A(n142), .ZN(n31) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n110), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n111), .A(n141), .ZN(n30) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n111), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n179), .B2(n103), .A(n140), .ZN(n3) );
  NAND2_X1 U21 ( .A1(data_in[29]), .A2(n110), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n153), .B2(n103), .A(n139), .ZN(n29) );
  NAND2_X1 U23 ( .A1(data_in[3]), .A2(n111), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n154), .B2(n103), .A(n138), .ZN(n28) );
  NAND2_X1 U25 ( .A1(data_in[4]), .A2(n111), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n155), .B2(ld), .A(n137), .ZN(n27) );
  NAND2_X1 U27 ( .A1(data_in[5]), .A2(n111), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n156), .B2(n110), .A(n136), .ZN(n26) );
  NAND2_X1 U29 ( .A1(data_in[6]), .A2(n111), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n157), .B2(n103), .A(n135), .ZN(n25) );
  NAND2_X1 U31 ( .A1(data_in[7]), .A2(n110), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n158), .B2(n103), .A(n134), .ZN(n24) );
  NAND2_X1 U33 ( .A1(data_in[8]), .A2(n111), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n159), .B2(n103), .A(n133), .ZN(n23) );
  NAND2_X1 U35 ( .A1(data_in[9]), .A2(n110), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n160), .B2(n103), .A(n132), .ZN(n22) );
  NAND2_X1 U37 ( .A1(data_in[10]), .A2(n110), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n161), .B2(n110), .A(n131), .ZN(n21) );
  NAND2_X1 U39 ( .A1(data_in[11]), .A2(n110), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n162), .B2(n111), .A(n130), .ZN(n20) );
  NAND2_X1 U41 ( .A1(data_in[12]), .A2(n110), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n180), .B2(n111), .A(n129), .ZN(n2) );
  NAND2_X1 U43 ( .A1(data_in[30]), .A2(n110), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n163), .B2(n110), .A(n128), .ZN(n19) );
  NAND2_X1 U45 ( .A1(data_in[13]), .A2(n110), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n164), .B2(n103), .A(n127), .ZN(n18) );
  NAND2_X1 U47 ( .A1(data_in[14]), .A2(n110), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n165), .B2(n110), .A(n126), .ZN(n17) );
  NAND2_X1 U49 ( .A1(data_in[15]), .A2(n111), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n166), .B2(n110), .A(n125), .ZN(n16) );
  NAND2_X1 U51 ( .A1(data_in[16]), .A2(n111), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n167), .B2(ld), .A(n124), .ZN(n15) );
  NAND2_X1 U53 ( .A1(data_in[17]), .A2(n110), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n168), .B2(n110), .A(n123), .ZN(n14) );
  NAND2_X1 U55 ( .A1(data_in[18]), .A2(n111), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n169), .B2(n111), .A(n122), .ZN(n13) );
  NAND2_X1 U57 ( .A1(data_in[19]), .A2(n111), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n170), .B2(n110), .A(n121), .ZN(n12) );
  NAND2_X1 U59 ( .A1(data_in[20]), .A2(n111), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n171), .B2(n103), .A(n120), .ZN(n11) );
  NAND2_X1 U61 ( .A1(data_in[21]), .A2(n111), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n172), .B2(ld), .A(n119), .ZN(n10) );
  NAND2_X1 U63 ( .A1(data_in[22]), .A2(n110), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n181), .B2(n103), .A(n118), .ZN(n1) );
  NAND2_X1 U65 ( .A1(data_in[31]), .A2(n110), .ZN(n118) );
  CLKBUF_X1 U69 ( .A(n111), .Z(n103) );
  CLKBUF_X1 U79 ( .A(rst), .Z(n116) );
  CLKBUF_X1 U80 ( .A(rst), .Z(n117) );
  CLKBUF_X1 U82 ( .A(ld), .Z(n110) );
  CLKBUF_X1 U83 ( .A(ld), .Z(n111) );
  DFFR_X1 \data_out_reg[29]  ( .D(n3), .CK(clk), .RN(n117), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n4), .CK(clk), .RN(n117), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n5), .CK(clk), .RN(n117), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n6), .CK(clk), .RN(n117), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n7), .CK(clk), .RN(n117), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n8), .CK(clk), .RN(n117), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n9), .CK(clk), .RN(n117), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n10), .CK(clk), .RN(n117), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n11), .CK(clk), .RN(n116), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n12), .CK(clk), .RN(n116), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n13), .CK(clk), .RN(n116), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n14), .CK(clk), .RN(n116), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n15), .CK(clk), .RN(n116), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n16), .CK(clk), .RN(n116), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n17), .CK(clk), .RN(n116), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n18), .CK(clk), .RN(n116), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n19), .CK(clk), .RN(n116), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n20), .CK(clk), .RN(n116), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n21), .CK(clk), .RN(n116), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n22), .CK(clk), .RN(n116), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n23), .CK(clk), .RN(n117), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n24), .CK(clk), .RN(n116), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n25), .CK(clk), .RN(n117), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n26), .CK(clk), .RN(n116), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n27), .CK(clk), .RN(n117), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n28), .CK(clk), .RN(n116), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n29), .CK(clk), .RN(n117), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n30), .CK(clk), .RN(n116), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n31), .CK(clk), .RN(n117), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n150) );
  DFFR_X1 \data_out_reg[31]  ( .D(n1), .CK(clk), .RN(n117), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n2), .CK(clk), .RN(n117), .Q(data_out[30]), 
        .QN(n180) );
endmodule


module cpsr ( clk, rst, ld, FL3, FL2, FL1, FL0, N, Z, C, V );
  input clk, rst, ld, FL3, FL2, FL1, FL0;
  output N, Z, C, V;
  wire   n9, n10, n11, n12, n1, n2, n3, n4, n5, n6, net83109, net83514, n7, n8,
         n13;

  OAI21_X1 U2 ( .B1(n4), .B2(ld), .A(n5), .ZN(n9) );
  NAND2_X1 U3 ( .A1(ld), .A2(FL1), .ZN(n5) );
  NAND2_X1 U5 ( .A1(FL0), .A2(ld), .ZN(n6) );
  NAND2_X1 U7 ( .A1(FL3), .A2(ld), .ZN(n7) );
  NAND2_X1 U9 ( .A1(FL2), .A2(ld), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n8), .A2(net83109), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n7), .A2(net83514), .ZN(n11) );
  OR2_X1 U8 ( .A1(n2), .A2(ld), .ZN(net83514) );
  OR2_X1 U10 ( .A1(n3), .A2(ld), .ZN(net83109) );
  OR2_X1 U11 ( .A1(n1), .A2(ld), .ZN(n13) );
  NAND2_X1 U12 ( .A1(n6), .A2(n13), .ZN(n12) );
  DFFR_X1 V_reg ( .D(n12), .CK(clk), .RN(rst), .Q(V), .QN(n1) );
  DFFR_X1 C_reg ( .D(n9), .CK(clk), .RN(rst), .Q(C), .QN(n4) );
  DFFR_X1 N_reg ( .D(n11), .CK(clk), .RN(rst), .Q(N), .QN(n2) );
  DFFR_X1 Z_reg ( .D(n10), .CK(clk), .RN(rst), .Q(Z), .QN(n3) );
endmodule


module gen_reg_N32_3 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n101, n102, n110, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  OAI21_X1 U2 ( .B1(n173), .B2(n101), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n102), .A2(data_in[23]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n174), .B2(ld), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[24]), .A2(n101), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n175), .B2(n101), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[25]), .A2(n101), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n176), .B2(n101), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[26]), .A2(n101), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n177), .B2(n101), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[27]), .A2(n102), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n178), .B2(n102), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[28]), .A2(n101), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n110), .A(n143), .ZN(n32) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n101), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n102), .A(n142), .ZN(n31) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n102), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n102), .A(n141), .ZN(n30) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n102), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n179), .B2(n110), .A(n140), .ZN(n3) );
  NAND2_X1 U21 ( .A1(data_in[29]), .A2(n102), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n153), .B2(n110), .A(n139), .ZN(n29) );
  NAND2_X1 U23 ( .A1(data_in[3]), .A2(n110), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n154), .B2(n102), .A(n138), .ZN(n28) );
  NAND2_X1 U25 ( .A1(data_in[4]), .A2(n101), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n155), .B2(n110), .A(n137), .ZN(n27) );
  NAND2_X1 U27 ( .A1(data_in[5]), .A2(n110), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n156), .B2(n102), .A(n136), .ZN(n26) );
  NAND2_X1 U29 ( .A1(data_in[6]), .A2(n101), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n157), .B2(n102), .A(n135), .ZN(n25) );
  NAND2_X1 U31 ( .A1(data_in[7]), .A2(n110), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n158), .B2(n102), .A(n134), .ZN(n24) );
  NAND2_X1 U33 ( .A1(data_in[8]), .A2(n110), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n159), .B2(n110), .A(n133), .ZN(n23) );
  NAND2_X1 U35 ( .A1(data_in[9]), .A2(n110), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n160), .B2(n101), .A(n132), .ZN(n22) );
  NAND2_X1 U37 ( .A1(data_in[10]), .A2(n102), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n161), .B2(n110), .A(n131), .ZN(n21) );
  NAND2_X1 U39 ( .A1(data_in[11]), .A2(n110), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n162), .B2(n102), .A(n130), .ZN(n20) );
  NAND2_X1 U41 ( .A1(data_in[12]), .A2(n110), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n180), .B2(n101), .A(n129), .ZN(n2) );
  NAND2_X1 U43 ( .A1(data_in[30]), .A2(n101), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n163), .B2(ld), .A(n128), .ZN(n19) );
  NAND2_X1 U45 ( .A1(data_in[13]), .A2(n101), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n164), .B2(n110), .A(n127), .ZN(n18) );
  NAND2_X1 U47 ( .A1(data_in[14]), .A2(n101), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n165), .B2(n101), .A(n126), .ZN(n17) );
  NAND2_X1 U49 ( .A1(data_in[15]), .A2(n102), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n166), .B2(n102), .A(n125), .ZN(n16) );
  NAND2_X1 U51 ( .A1(data_in[16]), .A2(n110), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n167), .B2(n102), .A(n124), .ZN(n15) );
  NAND2_X1 U53 ( .A1(data_in[17]), .A2(n102), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n168), .B2(n102), .A(n123), .ZN(n14) );
  NAND2_X1 U55 ( .A1(data_in[18]), .A2(ld), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n169), .B2(n102), .A(n122), .ZN(n13) );
  NAND2_X1 U57 ( .A1(data_in[19]), .A2(n102), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n170), .B2(n101), .A(n121), .ZN(n12) );
  NAND2_X1 U59 ( .A1(data_in[20]), .A2(n110), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n171), .B2(n101), .A(n120), .ZN(n11) );
  NAND2_X1 U61 ( .A1(data_in[21]), .A2(n101), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n172), .B2(n101), .A(n119), .ZN(n10) );
  NAND2_X1 U63 ( .A1(data_in[22]), .A2(n102), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n181), .B2(n101), .A(n118), .ZN(n1) );
  NAND2_X1 U65 ( .A1(data_in[31]), .A2(n110), .ZN(n118) );
  CLKBUF_X1 U68 ( .A(ld), .Z(n102) );
  CLKBUF_X1 U73 ( .A(ld), .Z(n101) );
  CLKBUF_X1 U79 ( .A(rst), .Z(n116) );
  CLKBUF_X1 U80 ( .A(rst), .Z(n117) );
  CLKBUF_X1 U82 ( .A(ld), .Z(n110) );
  DFFR_X1 \data_out_reg[31]  ( .D(n1), .CK(clk), .RN(n117), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n2), .CK(clk), .RN(n117), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n3), .CK(clk), .RN(n117), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n4), .CK(clk), .RN(n117), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n5), .CK(clk), .RN(n117), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n6), .CK(clk), .RN(n117), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n7), .CK(clk), .RN(n117), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n8), .CK(clk), .RN(n117), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n9), .CK(clk), .RN(n117), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n10), .CK(clk), .RN(n117), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n11), .CK(clk), .RN(n116), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n12), .CK(clk), .RN(n116), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n13), .CK(clk), .RN(n116), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n14), .CK(clk), .RN(n116), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n15), .CK(clk), .RN(n116), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n16), .CK(clk), .RN(n116), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n17), .CK(clk), .RN(n116), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n18), .CK(clk), .RN(n116), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n19), .CK(clk), .RN(n116), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n20), .CK(clk), .RN(n116), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n21), .CK(clk), .RN(n116), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n22), .CK(clk), .RN(n117), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n23), .CK(clk), .RN(n116), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n24), .CK(clk), .RN(n117), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n25), .CK(clk), .RN(n116), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n26), .CK(clk), .RN(n117), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n27), .CK(clk), .RN(n116), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n28), .CK(clk), .RN(n117), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n29), .CK(clk), .RN(n116), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n30), .CK(clk), .RN(n117), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n31), .CK(clk), .RN(n116), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n32), .CK(clk), .RN(n117), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N5_2 ( clk, rst, ld, data_in, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26;

  OAI21_X1 U2 ( .B1(n22), .B2(n16), .A(n21), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n16), .A2(data_in[0]), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n23), .B2(n16), .A(n20), .ZN(n4) );
  NAND2_X1 U5 ( .A1(data_in[1]), .A2(n16), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(n16), .A(n19), .ZN(n3) );
  NAND2_X1 U7 ( .A1(data_in[2]), .A2(n16), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n25), .B2(n16), .A(n18), .ZN(n2) );
  NAND2_X1 U9 ( .A1(data_in[3]), .A2(n16), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n26), .B2(n16), .A(n17), .ZN(n1) );
  NAND2_X1 U11 ( .A1(data_in[4]), .A2(n16), .ZN(n17) );
  CLKBUF_X1 U12 ( .A(ld), .Z(n16) );
  DFFR_X1 \data_out_reg[4]  ( .D(n1), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n26) );
  DFFR_X1 \data_out_reg[3]  ( .D(n2), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n25) );
  DFFR_X1 \data_out_reg[2]  ( .D(n3), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n24) );
  DFFR_X1 \data_out_reg[1]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n23) );
  DFFR_X1 \data_out_reg[0]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n22) );
endmodule


module gen_mux21_N32_1 ( sel, x, y, m );
  input [31:0] x;
  input [31:0] y;
  output [31:0] m;
  input sel;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, net74348, net74349, net75107, net75105, net75111, net76798,
         net76797, net76802, net76801, net76806, net110268, n33, n41, n42, n66
;
  assign m[30] = net74348;
  assign m[31] = net74349;
  assign net75111 = sel;

  AOI22_X1 U34 ( .A1(x[9]), .A2(net76806), .B1(y[9]), .B2(net75111), .ZN(n34)
         );
  AOI22_X1 U35 ( .A1(x[8]), .A2(net76806), .B1(y[8]), .B2(net75111), .ZN(n35)
         );
  AOI22_X1 U36 ( .A1(x[7]), .A2(net76806), .B1(y[7]), .B2(net75111), .ZN(n36)
         );
  AOI22_X1 U37 ( .A1(x[6]), .A2(net76806), .B1(y[6]), .B2(net75111), .ZN(n37)
         );
  AOI22_X1 U38 ( .A1(x[5]), .A2(net76806), .B1(y[5]), .B2(net75111), .ZN(n38)
         );
  AOI22_X1 U39 ( .A1(x[4]), .A2(net76806), .B1(y[4]), .B2(net75111), .ZN(n39)
         );
  AOI22_X1 U40 ( .A1(x[3]), .A2(net76806), .B1(y[3]), .B2(net75111), .ZN(n40)
         );
  AOI22_X1 U43 ( .A1(x[2]), .A2(net76806), .B1(y[2]), .B2(net75111), .ZN(n43)
         );
  AOI22_X1 U44 ( .A1(x[29]), .A2(net76806), .B1(y[29]), .B2(net75111), .ZN(n44) );
  AOI22_X1 U45 ( .A1(x[28]), .A2(net76801), .B1(y[28]), .B2(net75111), .ZN(n45) );
  AOI22_X1 U46 ( .A1(x[27]), .A2(net76802), .B1(y[27]), .B2(net75111), .ZN(n46) );
  AOI22_X1 U47 ( .A1(x[26]), .A2(net76801), .B1(y[26]), .B2(net75111), .ZN(n47) );
  AOI22_X1 U48 ( .A1(x[25]), .A2(net76802), .B1(y[25]), .B2(net75111), .ZN(n48) );
  AOI22_X1 U49 ( .A1(x[24]), .A2(net76801), .B1(y[24]), .B2(net75111), .ZN(n49) );
  AOI22_X1 U50 ( .A1(x[23]), .A2(net76802), .B1(y[23]), .B2(net75111), .ZN(n50) );
  AOI22_X1 U51 ( .A1(x[22]), .A2(net76801), .B1(y[22]), .B2(net75111), .ZN(n51) );
  AOI22_X1 U52 ( .A1(x[21]), .A2(net76802), .B1(y[21]), .B2(net75105), .ZN(n52) );
  AOI22_X1 U53 ( .A1(x[20]), .A2(net76801), .B1(y[20]), .B2(net75105), .ZN(n53) );
  AOI22_X1 U54 ( .A1(x[1]), .A2(net76802), .B1(y[1]), .B2(net75105), .ZN(n54)
         );
  AOI22_X1 U55 ( .A1(x[19]), .A2(net76801), .B1(y[19]), .B2(net75105), .ZN(n55) );
  AOI22_X1 U56 ( .A1(x[18]), .A2(net76798), .B1(y[18]), .B2(net75105), .ZN(n56) );
  AOI22_X1 U57 ( .A1(x[17]), .A2(net76797), .B1(y[17]), .B2(net75105), .ZN(n57) );
  AOI22_X1 U58 ( .A1(x[16]), .A2(net76798), .B1(y[16]), .B2(net75105), .ZN(n58) );
  AOI22_X1 U59 ( .A1(x[15]), .A2(net76797), .B1(y[15]), .B2(net75107), .ZN(n59) );
  AOI22_X1 U60 ( .A1(x[14]), .A2(net76798), .B1(y[14]), .B2(net75107), .ZN(n60) );
  AOI22_X1 U61 ( .A1(x[13]), .A2(net76797), .B1(y[13]), .B2(net75107), .ZN(n61) );
  AOI22_X1 U62 ( .A1(x[12]), .A2(net76798), .B1(y[12]), .B2(net75107), .ZN(n62) );
  AOI22_X1 U63 ( .A1(x[11]), .A2(net76797), .B1(y[11]), .B2(net75107), .ZN(n63) );
  AOI22_X1 U64 ( .A1(x[10]), .A2(net76798), .B1(y[10]), .B2(net75107), .ZN(n64) );
  AOI22_X1 U65 ( .A1(x[0]), .A2(net76797), .B1(y[0]), .B2(net75107), .ZN(n65)
         );
  NAND2_X1 U1 ( .A1(y[30]), .A2(net75105), .ZN(n33) );
  NAND2_X1 U2 ( .A1(n33), .A2(n41), .ZN(net74348) );
  NAND2_X1 U5 ( .A1(x[30]), .A2(net110268), .ZN(n41) );
  NAND2_X1 U6 ( .A1(n42), .A2(n66), .ZN(net74349) );
  NAND2_X1 U7 ( .A1(x[31]), .A2(net110268), .ZN(n66) );
  INV_X1 U8 ( .A(net75111), .ZN(net110268) );
  NAND2_X1 U10 ( .A1(y[31]), .A2(net75107), .ZN(n42) );
  CLKBUF_X1 U12 ( .A(net110268), .Z(net76801) );
  CLKBUF_X1 U13 ( .A(net110268), .Z(net76797) );
  CLKBUF_X1 U14 ( .A(net110268), .Z(net76798) );
  CLKBUF_X1 U15 ( .A(net110268), .Z(net76802) );
  CLKBUF_X1 U16 ( .A(net75111), .Z(net75107) );
  CLKBUF_X1 U17 ( .A(net75111), .Z(net75105) );
  INV_X1 U18 ( .A(n44), .ZN(m[29]) );
  INV_X1 U19 ( .A(n45), .ZN(m[28]) );
  INV_X1 U20 ( .A(n46), .ZN(m[27]) );
  INV_X1 U21 ( .A(n47), .ZN(m[26]) );
  INV_X1 U22 ( .A(n48), .ZN(m[25]) );
  INV_X1 U23 ( .A(n49), .ZN(m[24]) );
  INV_X1 U24 ( .A(n50), .ZN(m[23]) );
  INV_X1 U25 ( .A(n51), .ZN(m[22]) );
  INV_X1 U26 ( .A(n52), .ZN(m[21]) );
  INV_X1 U27 ( .A(n53), .ZN(m[20]) );
  INV_X1 U28 ( .A(n60), .ZN(m[14]) );
  INV_X1 U29 ( .A(n59), .ZN(m[15]) );
  INV_X1 U30 ( .A(n58), .ZN(m[16]) );
  INV_X1 U31 ( .A(n55), .ZN(m[19]) );
  INV_X1 U32 ( .A(n56), .ZN(m[18]) );
  INV_X1 U33 ( .A(n57), .ZN(m[17]) );
  INV_X1 U41 ( .A(n65), .ZN(m[0]) );
  INV_X1 U42 ( .A(n35), .ZN(m[8]) );
  INV_X1 U66 ( .A(n34), .ZN(m[9]) );
  INV_X1 U67 ( .A(n64), .ZN(m[10]) );
  INV_X1 U68 ( .A(n63), .ZN(m[11]) );
  INV_X1 U69 ( .A(n62), .ZN(m[12]) );
  INV_X1 U70 ( .A(n61), .ZN(m[13]) );
  INV_X1 U71 ( .A(n39), .ZN(m[4]) );
  INV_X1 U72 ( .A(n38), .ZN(m[5]) );
  INV_X1 U73 ( .A(n37), .ZN(m[6]) );
  INV_X1 U74 ( .A(n36), .ZN(m[7]) );
  INV_X1 U75 ( .A(n54), .ZN(m[1]) );
  INV_X1 U76 ( .A(n43), .ZN(m[2]) );
  INV_X1 U77 ( .A(n40), .ZN(m[3]) );
  INV_X1 U3 ( .A(net75111), .ZN(net76806) );
endmodule


module EXE_STAGE_N_BITS_DATA32_RF_ADDR5 ( CLK, RST, MUXA_SEL, MUXB_SEL, 
        EXE_OUTREG_EN, EQ_COND, JUMP_EN, .ALU_OPCODE({\ALU_OPCODE[6] , 
        \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , 
        \ALU_OPCODE[1] , \ALU_OPCODE[0] }), NPC2_IN, NPC1_MUXA_IN, 
        REGA_MUXA_IN, REGB_MUXB_IN, IMM_MUXB_IN, PAD_IN, IR2_IN, JUMP_MUX_IN_0, 
        NPC2_OUT, ALU_OUT, PAD_OUT, IR2_OUT, ADDR_MUX_OUT, N_FLAG, Z_FLAG, 
        C_FLAG, V_FLAG );
  input [31:0] NPC2_IN;
  input [31:0] NPC1_MUXA_IN;
  input [31:0] REGA_MUXA_IN;
  input [31:0] REGB_MUXB_IN;
  input [31:0] IMM_MUXB_IN;
  input [31:0] PAD_IN;
  input [4:0] IR2_IN;
  input [31:0] JUMP_MUX_IN_0;
  output [31:0] NPC2_OUT;
  output [31:0] ALU_OUT;
  output [31:0] PAD_OUT;
  output [4:0] IR2_OUT;
  output [31:0] ADDR_MUX_OUT;
  input CLK, RST, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN,
         \ALU_OPCODE[6] , \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] ;
  output N_FLAG, Z_FLAG, C_FLAG, V_FLAG;
  wire   BRANCH_TAKEN, COND_OUT, NEG_INT, ZERO_INT, CARRY_INT, OVF_INT;
  wire   [6:0] ALU_OPCODE;
  wire   [31:0] MUXA_OUT_INT;
  wire   [31:0] MUXB_OUT_INT;
  wire   [31:0] ALU_OUT_INT;

  gen_reg_N32_5 NPC2 ( .clk(CLK), .rst(RST), .ld(EXE_OUTREG_EN), .data_in(
        NPC2_IN), .data_out(NPC2_OUT) );
  zero_check_N32 ZERO ( .data_in(REGA_MUXA_IN), .ctrl_out(BRANCH_TAKEN) );
  cond_branch COND ( .cond_in(EQ_COND), .jump_in(JUMP_EN), .ctrl_in(
        BRANCH_TAKEN), .ctrl_out(COND_OUT) );
  gen_mux21_N32_0 MUXA ( .sel(MUXA_SEL), .x(NPC1_MUXA_IN), .y(REGA_MUXA_IN), 
        .m(MUXA_OUT_INT) );
  gen_mux21_N32_2 MUXB ( .sel(MUXB_SEL), .x(REGB_MUXB_IN), .y(IMM_MUXB_IN), 
        .m(MUXB_OUT_INT) );
  ALU_N32 ALRITH_LOG_U ( .ALU_OPCODE({\ALU_OPCODE[6] , \ALU_OPCODE[5] , 
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), .DATA1(MUXA_OUT_INT), .DATA2(MUXB_OUT_INT), .NEG(
        NEG_INT), .ZERO(ZERO_INT), .CARRY(CARRY_INT), .OVF(OVF_INT), .OUTALU(
        ALU_OUT_INT) );
  gen_reg_N32_4 ALU_OUTPUT ( .clk(CLK), .rst(RST), .ld(EXE_OUTREG_EN), 
        .data_in(ALU_OUT_INT), .data_out(ALU_OUT) );
  cpsr ALU_FLAGS ( .clk(CLK), .rst(RST), .ld(EXE_OUTREG_EN), .FL3(NEG_INT), 
        .FL2(ZERO_INT), .FL1(CARRY_INT), .FL0(OVF_INT), .N(N_FLAG), .Z(Z_FLAG), 
        .C(C_FLAG), .V(V_FLAG) );
  gen_reg_N32_3 PAD ( .clk(CLK), .rst(RST), .ld(EXE_OUTREG_EN), .data_in(
        PAD_IN), .data_out(PAD_OUT) );
  gen_reg_N5_2 IR2 ( .clk(CLK), .rst(RST), .ld(EXE_OUTREG_EN), .data_in(IR2_IN), .data_out(IR2_OUT) );
  gen_mux21_N32_1 ADDR_MUX ( .sel(COND_OUT), .x(JUMP_MUX_IN_0), .y(ALU_OUT_INT), .m(ADDR_MUX_OUT) );
endmodule


module gen_reg_N32_2 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n99, n100, n109, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181;

  OAI21_X1 U2 ( .B1(n173), .B2(n109), .A(n149), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n100), .A2(data_in[23]), .ZN(n149) );
  OAI21_X1 U4 ( .B1(n174), .B2(ld), .A(n148), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[24]), .A2(n109), .ZN(n148) );
  OAI21_X1 U6 ( .B1(n175), .B2(n99), .A(n147), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[25]), .A2(n109), .ZN(n147) );
  OAI21_X1 U8 ( .B1(n176), .B2(n109), .A(n146), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[26]), .A2(n109), .ZN(n146) );
  OAI21_X1 U10 ( .B1(n177), .B2(n99), .A(n145), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[27]), .A2(n99), .ZN(n145) );
  OAI21_X1 U12 ( .B1(n178), .B2(n109), .A(n144), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[28]), .A2(n99), .ZN(n144) );
  OAI21_X1 U14 ( .B1(n150), .B2(n100), .A(n143), .ZN(n32) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(n99), .ZN(n143) );
  OAI21_X1 U16 ( .B1(n151), .B2(n100), .A(n142), .ZN(n31) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(n99), .ZN(n142) );
  OAI21_X1 U18 ( .B1(n152), .B2(n109), .A(n141), .ZN(n30) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(n99), .ZN(n141) );
  OAI21_X1 U20 ( .B1(n179), .B2(n100), .A(n140), .ZN(n3) );
  NAND2_X1 U21 ( .A1(data_in[29]), .A2(n99), .ZN(n140) );
  OAI21_X1 U22 ( .B1(n153), .B2(n100), .A(n139), .ZN(n29) );
  NAND2_X1 U23 ( .A1(data_in[3]), .A2(n100), .ZN(n139) );
  OAI21_X1 U24 ( .B1(n154), .B2(n109), .A(n138), .ZN(n28) );
  NAND2_X1 U25 ( .A1(data_in[4]), .A2(n99), .ZN(n138) );
  OAI21_X1 U26 ( .B1(n155), .B2(n99), .A(n137), .ZN(n27) );
  NAND2_X1 U27 ( .A1(data_in[5]), .A2(n100), .ZN(n137) );
  OAI21_X1 U28 ( .B1(n156), .B2(n99), .A(n136), .ZN(n26) );
  NAND2_X1 U29 ( .A1(data_in[6]), .A2(n99), .ZN(n136) );
  OAI21_X1 U30 ( .B1(n157), .B2(n100), .A(n135), .ZN(n25) );
  NAND2_X1 U31 ( .A1(data_in[7]), .A2(n100), .ZN(n135) );
  OAI21_X1 U32 ( .B1(n158), .B2(n100), .A(n134), .ZN(n24) );
  NAND2_X1 U33 ( .A1(data_in[8]), .A2(n99), .ZN(n134) );
  OAI21_X1 U34 ( .B1(n159), .B2(n100), .A(n133), .ZN(n23) );
  NAND2_X1 U35 ( .A1(data_in[9]), .A2(n100), .ZN(n133) );
  OAI21_X1 U36 ( .B1(n160), .B2(n100), .A(n132), .ZN(n22) );
  NAND2_X1 U37 ( .A1(data_in[10]), .A2(n99), .ZN(n132) );
  OAI21_X1 U38 ( .B1(n161), .B2(n109), .A(n131), .ZN(n21) );
  NAND2_X1 U39 ( .A1(data_in[11]), .A2(n100), .ZN(n131) );
  OAI21_X1 U40 ( .B1(n162), .B2(n100), .A(n130), .ZN(n20) );
  NAND2_X1 U41 ( .A1(data_in[12]), .A2(n99), .ZN(n130) );
  OAI21_X1 U42 ( .B1(n180), .B2(n99), .A(n129), .ZN(n2) );
  NAND2_X1 U43 ( .A1(data_in[30]), .A2(n109), .ZN(n129) );
  OAI21_X1 U44 ( .B1(n163), .B2(n100), .A(n128), .ZN(n19) );
  NAND2_X1 U45 ( .A1(data_in[13]), .A2(n109), .ZN(n128) );
  OAI21_X1 U46 ( .B1(n164), .B2(n99), .A(n127), .ZN(n18) );
  NAND2_X1 U47 ( .A1(data_in[14]), .A2(n109), .ZN(n127) );
  OAI21_X1 U48 ( .B1(n165), .B2(n109), .A(n126), .ZN(n17) );
  NAND2_X1 U49 ( .A1(data_in[15]), .A2(n109), .ZN(n126) );
  OAI21_X1 U50 ( .B1(n166), .B2(n100), .A(n125), .ZN(n16) );
  NAND2_X1 U51 ( .A1(data_in[16]), .A2(n99), .ZN(n125) );
  OAI21_X1 U52 ( .B1(n167), .B2(n99), .A(n124), .ZN(n15) );
  NAND2_X1 U53 ( .A1(data_in[17]), .A2(n109), .ZN(n124) );
  OAI21_X1 U54 ( .B1(n168), .B2(n100), .A(n123), .ZN(n14) );
  NAND2_X1 U55 ( .A1(data_in[18]), .A2(n100), .ZN(n123) );
  OAI21_X1 U56 ( .B1(n169), .B2(n99), .A(n122), .ZN(n13) );
  NAND2_X1 U57 ( .A1(data_in[19]), .A2(n109), .ZN(n122) );
  OAI21_X1 U58 ( .B1(n170), .B2(n100), .A(n121), .ZN(n12) );
  NAND2_X1 U59 ( .A1(data_in[20]), .A2(n100), .ZN(n121) );
  OAI21_X1 U60 ( .B1(n171), .B2(n100), .A(n120), .ZN(n11) );
  NAND2_X1 U61 ( .A1(data_in[21]), .A2(n109), .ZN(n120) );
  OAI21_X1 U62 ( .B1(n172), .B2(n99), .A(n119), .ZN(n10) );
  NAND2_X1 U63 ( .A1(data_in[22]), .A2(n99), .ZN(n119) );
  OAI21_X1 U64 ( .B1(n181), .B2(n100), .A(n118), .ZN(n1) );
  NAND2_X1 U65 ( .A1(data_in[31]), .A2(n99), .ZN(n118) );
  CLKBUF_X1 U70 ( .A(ld), .Z(n99) );
  CLKBUF_X1 U74 ( .A(ld), .Z(n100) );
  CLKBUF_X1 U81 ( .A(ld), .Z(n109) );
  DFFR_X1 \data_out_reg[31]  ( .D(n1), .CK(clk), .RN(rst), .Q(data_out[31]), 
        .QN(n181) );
  DFFR_X1 \data_out_reg[30]  ( .D(n2), .CK(clk), .RN(rst), .Q(data_out[30]), 
        .QN(n180) );
  DFFR_X1 \data_out_reg[29]  ( .D(n3), .CK(clk), .RN(rst), .Q(data_out[29]), 
        .QN(n179) );
  DFFR_X1 \data_out_reg[28]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[28]), 
        .QN(n178) );
  DFFR_X1 \data_out_reg[27]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[27]), 
        .QN(n177) );
  DFFR_X1 \data_out_reg[26]  ( .D(n6), .CK(clk), .RN(rst), .Q(data_out[26]), 
        .QN(n176) );
  DFFR_X1 \data_out_reg[25]  ( .D(n7), .CK(clk), .RN(rst), .Q(data_out[25]), 
        .QN(n175) );
  DFFR_X1 \data_out_reg[24]  ( .D(n8), .CK(clk), .RN(rst), .Q(data_out[24]), 
        .QN(n174) );
  DFFR_X1 \data_out_reg[23]  ( .D(n9), .CK(clk), .RN(rst), .Q(data_out[23]), 
        .QN(n173) );
  DFFR_X1 \data_out_reg[22]  ( .D(n10), .CK(clk), .RN(rst), .Q(data_out[22]), 
        .QN(n172) );
  DFFR_X1 \data_out_reg[21]  ( .D(n11), .CK(clk), .RN(rst), .Q(data_out[21]), 
        .QN(n171) );
  DFFR_X1 \data_out_reg[20]  ( .D(n12), .CK(clk), .RN(rst), .Q(data_out[20]), 
        .QN(n170) );
  DFFR_X1 \data_out_reg[19]  ( .D(n13), .CK(clk), .RN(rst), .Q(data_out[19]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[18]  ( .D(n14), .CK(clk), .RN(rst), .Q(data_out[18]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[17]  ( .D(n15), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[16]  ( .D(n16), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[15]  ( .D(n17), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[14]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[13]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[12]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[12]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[11]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[11]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[10]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[10]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[9]  ( .D(n23), .CK(clk), .RN(rst), .Q(data_out[9]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[8]  ( .D(n24), .CK(clk), .RN(rst), .Q(data_out[8]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[7]  ( .D(n25), .CK(clk), .RN(rst), .Q(data_out[7]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[6]  ( .D(n26), .CK(clk), .RN(rst), .Q(data_out[6]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[5]  ( .D(n27), .CK(clk), .RN(rst), .Q(data_out[5]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[4]  ( .D(n28), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[3]  ( .D(n29), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[2]  ( .D(n30), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[1]  ( .D(n31), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[0]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n150) );
endmodule


module gen_reg_N32_1 ( clk, rst, ld, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n101, n102, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169;

  OAI21_X1 U2 ( .B1(n161), .B2(n102), .A(n137), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n101), .A2(data_in[23]), .ZN(n137) );
  OAI21_X1 U4 ( .B1(n162), .B2(n102), .A(n136), .ZN(n8) );
  NAND2_X1 U5 ( .A1(data_in[24]), .A2(n102), .ZN(n136) );
  OAI21_X1 U6 ( .B1(n163), .B2(n102), .A(n135), .ZN(n7) );
  NAND2_X1 U7 ( .A1(data_in[25]), .A2(ld), .ZN(n135) );
  OAI21_X1 U8 ( .B1(n164), .B2(n102), .A(n134), .ZN(n6) );
  NAND2_X1 U9 ( .A1(data_in[26]), .A2(n101), .ZN(n134) );
  OAI21_X1 U10 ( .B1(n165), .B2(n101), .A(n133), .ZN(n5) );
  NAND2_X1 U11 ( .A1(data_in[27]), .A2(n102), .ZN(n133) );
  OAI21_X1 U12 ( .B1(n166), .B2(n101), .A(n132), .ZN(n4) );
  NAND2_X1 U13 ( .A1(data_in[28]), .A2(ld), .ZN(n132) );
  OAI21_X1 U14 ( .B1(n138), .B2(n101), .A(n131), .ZN(n32) );
  NAND2_X1 U15 ( .A1(data_in[0]), .A2(ld), .ZN(n131) );
  OAI21_X1 U16 ( .B1(n139), .B2(n101), .A(n130), .ZN(n31) );
  NAND2_X1 U17 ( .A1(data_in[1]), .A2(ld), .ZN(n130) );
  OAI21_X1 U18 ( .B1(n140), .B2(n102), .A(n129), .ZN(n30) );
  NAND2_X1 U19 ( .A1(data_in[2]), .A2(ld), .ZN(n129) );
  OAI21_X1 U20 ( .B1(n167), .B2(n101), .A(n128), .ZN(n3) );
  NAND2_X1 U21 ( .A1(data_in[29]), .A2(n102), .ZN(n128) );
  OAI21_X1 U22 ( .B1(n141), .B2(n102), .A(n127), .ZN(n29) );
  NAND2_X1 U23 ( .A1(data_in[3]), .A2(ld), .ZN(n127) );
  OAI21_X1 U24 ( .B1(n142), .B2(n102), .A(n126), .ZN(n28) );
  NAND2_X1 U25 ( .A1(data_in[4]), .A2(ld), .ZN(n126) );
  OAI21_X1 U26 ( .B1(n143), .B2(n101), .A(n125), .ZN(n27) );
  NAND2_X1 U27 ( .A1(data_in[5]), .A2(ld), .ZN(n125) );
  OAI21_X1 U28 ( .B1(n144), .B2(n102), .A(n124), .ZN(n26) );
  NAND2_X1 U29 ( .A1(data_in[6]), .A2(ld), .ZN(n124) );
  OAI21_X1 U30 ( .B1(n145), .B2(n101), .A(n123), .ZN(n25) );
  NAND2_X1 U31 ( .A1(data_in[7]), .A2(ld), .ZN(n123) );
  OAI21_X1 U32 ( .B1(n146), .B2(n102), .A(n122), .ZN(n24) );
  NAND2_X1 U33 ( .A1(data_in[8]), .A2(ld), .ZN(n122) );
  OAI21_X1 U34 ( .B1(n147), .B2(n101), .A(n121), .ZN(n23) );
  NAND2_X1 U35 ( .A1(data_in[9]), .A2(ld), .ZN(n121) );
  OAI21_X1 U36 ( .B1(n148), .B2(n102), .A(n120), .ZN(n22) );
  NAND2_X1 U37 ( .A1(data_in[10]), .A2(ld), .ZN(n120) );
  OAI21_X1 U38 ( .B1(n149), .B2(n101), .A(n119), .ZN(n21) );
  NAND2_X1 U39 ( .A1(data_in[11]), .A2(n101), .ZN(n119) );
  OAI21_X1 U40 ( .B1(n150), .B2(n102), .A(n118), .ZN(n20) );
  NAND2_X1 U41 ( .A1(data_in[12]), .A2(n101), .ZN(n118) );
  OAI21_X1 U42 ( .B1(n168), .B2(n101), .A(n117), .ZN(n2) );
  NAND2_X1 U43 ( .A1(data_in[30]), .A2(ld), .ZN(n117) );
  OAI21_X1 U44 ( .B1(n151), .B2(n101), .A(n116), .ZN(n19) );
  NAND2_X1 U45 ( .A1(data_in[13]), .A2(ld), .ZN(n116) );
  OAI21_X1 U46 ( .B1(n152), .B2(n101), .A(n115), .ZN(n18) );
  NAND2_X1 U47 ( .A1(data_in[14]), .A2(n102), .ZN(n115) );
  OAI21_X1 U48 ( .B1(n153), .B2(n101), .A(n114), .ZN(n17) );
  NAND2_X1 U49 ( .A1(data_in[15]), .A2(n102), .ZN(n114) );
  OAI21_X1 U50 ( .B1(n154), .B2(n101), .A(n113), .ZN(n16) );
  NAND2_X1 U51 ( .A1(data_in[16]), .A2(n101), .ZN(n113) );
  OAI21_X1 U52 ( .B1(n155), .B2(n101), .A(n112), .ZN(n15) );
  NAND2_X1 U53 ( .A1(data_in[17]), .A2(n102), .ZN(n112) );
  OAI21_X1 U54 ( .B1(n156), .B2(n101), .A(n111), .ZN(n14) );
  NAND2_X1 U55 ( .A1(data_in[18]), .A2(n102), .ZN(n111) );
  OAI21_X1 U56 ( .B1(n157), .B2(n102), .A(n110), .ZN(n13) );
  NAND2_X1 U57 ( .A1(data_in[19]), .A2(ld), .ZN(n110) );
  OAI21_X1 U58 ( .B1(n158), .B2(n102), .A(n109), .ZN(n12) );
  NAND2_X1 U59 ( .A1(data_in[20]), .A2(ld), .ZN(n109) );
  OAI21_X1 U60 ( .B1(n159), .B2(n102), .A(n108), .ZN(n11) );
  NAND2_X1 U61 ( .A1(data_in[21]), .A2(ld), .ZN(n108) );
  OAI21_X1 U62 ( .B1(n160), .B2(n102), .A(n107), .ZN(n10) );
  NAND2_X1 U63 ( .A1(data_in[22]), .A2(ld), .ZN(n107) );
  OAI21_X1 U64 ( .B1(n169), .B2(n102), .A(n106), .ZN(n1) );
  NAND2_X1 U65 ( .A1(data_in[31]), .A2(n101), .ZN(n106) );
  CLKBUF_X1 U73 ( .A(ld), .Z(n101) );
  CLKBUF_X1 U74 ( .A(ld), .Z(n102) );
  DFFR_X1 \data_out_reg[31]  ( .D(n1), .CK(clk), .RN(rst), .Q(data_out[31]), 
        .QN(n169) );
  DFFR_X1 \data_out_reg[30]  ( .D(n2), .CK(clk), .RN(rst), .Q(data_out[30]), 
        .QN(n168) );
  DFFR_X1 \data_out_reg[29]  ( .D(n3), .CK(clk), .RN(rst), .Q(data_out[29]), 
        .QN(n167) );
  DFFR_X1 \data_out_reg[28]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[28]), 
        .QN(n166) );
  DFFR_X1 \data_out_reg[27]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[27]), 
        .QN(n165) );
  DFFR_X1 \data_out_reg[26]  ( .D(n6), .CK(clk), .RN(rst), .Q(data_out[26]), 
        .QN(n164) );
  DFFR_X1 \data_out_reg[25]  ( .D(n7), .CK(clk), .RN(rst), .Q(data_out[25]), 
        .QN(n163) );
  DFFR_X1 \data_out_reg[24]  ( .D(n8), .CK(clk), .RN(rst), .Q(data_out[24]), 
        .QN(n162) );
  DFFR_X1 \data_out_reg[23]  ( .D(n9), .CK(clk), .RN(rst), .Q(data_out[23]), 
        .QN(n161) );
  DFFR_X1 \data_out_reg[22]  ( .D(n10), .CK(clk), .RN(rst), .Q(data_out[22]), 
        .QN(n160) );
  DFFR_X1 \data_out_reg[21]  ( .D(n11), .CK(clk), .RN(rst), .Q(data_out[21]), 
        .QN(n159) );
  DFFR_X1 \data_out_reg[20]  ( .D(n12), .CK(clk), .RN(rst), .Q(data_out[20]), 
        .QN(n158) );
  DFFR_X1 \data_out_reg[19]  ( .D(n13), .CK(clk), .RN(rst), .Q(data_out[19]), 
        .QN(n157) );
  DFFR_X1 \data_out_reg[18]  ( .D(n14), .CK(clk), .RN(rst), .Q(data_out[18]), 
        .QN(n156) );
  DFFR_X1 \data_out_reg[17]  ( .D(n15), .CK(clk), .RN(rst), .Q(data_out[17]), 
        .QN(n155) );
  DFFR_X1 \data_out_reg[16]  ( .D(n16), .CK(clk), .RN(rst), .Q(data_out[16]), 
        .QN(n154) );
  DFFR_X1 \data_out_reg[15]  ( .D(n17), .CK(clk), .RN(rst), .Q(data_out[15]), 
        .QN(n153) );
  DFFR_X1 \data_out_reg[14]  ( .D(n18), .CK(clk), .RN(rst), .Q(data_out[14]), 
        .QN(n152) );
  DFFR_X1 \data_out_reg[13]  ( .D(n19), .CK(clk), .RN(rst), .Q(data_out[13]), 
        .QN(n151) );
  DFFR_X1 \data_out_reg[12]  ( .D(n20), .CK(clk), .RN(rst), .Q(data_out[12]), 
        .QN(n150) );
  DFFR_X1 \data_out_reg[11]  ( .D(n21), .CK(clk), .RN(rst), .Q(data_out[11]), 
        .QN(n149) );
  DFFR_X1 \data_out_reg[10]  ( .D(n22), .CK(clk), .RN(rst), .Q(data_out[10]), 
        .QN(n148) );
  DFFR_X1 \data_out_reg[9]  ( .D(n23), .CK(clk), .RN(rst), .Q(data_out[9]), 
        .QN(n147) );
  DFFR_X1 \data_out_reg[8]  ( .D(n24), .CK(clk), .RN(rst), .Q(data_out[8]), 
        .QN(n146) );
  DFFR_X1 \data_out_reg[7]  ( .D(n25), .CK(clk), .RN(rst), .Q(data_out[7]), 
        .QN(n145) );
  DFFR_X1 \data_out_reg[6]  ( .D(n26), .CK(clk), .RN(rst), .Q(data_out[6]), 
        .QN(n144) );
  DFFR_X1 \data_out_reg[5]  ( .D(n27), .CK(clk), .RN(rst), .Q(data_out[5]), 
        .QN(n143) );
  DFFR_X1 \data_out_reg[4]  ( .D(n28), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n142) );
  DFFR_X1 \data_out_reg[3]  ( .D(n29), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n141) );
  DFFR_X1 \data_out_reg[2]  ( .D(n30), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n140) );
  DFFR_X1 \data_out_reg[1]  ( .D(n31), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n139) );
  DFFR_X1 \data_out_reg[0]  ( .D(n32), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n138) );
endmodule


module gen_reg_N5_1 ( clk, rst, ld, data_in, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, rst, ld;
  wire   n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26;

  OAI21_X1 U2 ( .B1(n22), .B2(n16), .A(n21), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n16), .A2(data_in[0]), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n23), .B2(n16), .A(n20), .ZN(n4) );
  NAND2_X1 U5 ( .A1(data_in[1]), .A2(n16), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(n16), .A(n19), .ZN(n3) );
  NAND2_X1 U7 ( .A1(data_in[2]), .A2(n16), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n25), .B2(n16), .A(n18), .ZN(n2) );
  NAND2_X1 U9 ( .A1(data_in[3]), .A2(n16), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n26), .B2(n16), .A(n17), .ZN(n1) );
  NAND2_X1 U11 ( .A1(data_in[4]), .A2(n16), .ZN(n17) );
  CLKBUF_X1 U12 ( .A(ld), .Z(n16) );
  DFFR_X1 \data_out_reg[4]  ( .D(n1), .CK(clk), .RN(rst), .Q(data_out[4]), 
        .QN(n26) );
  DFFR_X1 \data_out_reg[3]  ( .D(n2), .CK(clk), .RN(rst), .Q(data_out[3]), 
        .QN(n25) );
  DFFR_X1 \data_out_reg[2]  ( .D(n3), .CK(clk), .RN(rst), .Q(data_out[2]), 
        .QN(n24) );
  DFFR_X1 \data_out_reg[1]  ( .D(n4), .CK(clk), .RN(rst), .Q(data_out[1]), 
        .QN(n23) );
  DFFR_X1 \data_out_reg[0]  ( .D(n5), .CK(clk), .RN(rst), .Q(data_out[0]), 
        .QN(n22) );
endmodule


module MEM_STAGE_N_BITS_DATA32_RF_ADDR5 ( CLK, RST, MEM_OUTREG_EN, BYTE_LEN_IN, 
        DRAM_WE, DRAM_WE_OUT, BYTE_LEN_OUT, ALU_OUTPUT_IN, MEM_DATA_IN, 
        MEM_DATA_OUT_INT, NPC_IN, IR_IN, IR_OUT, NPC_OUT, MEM_ADDR_OUT, 
        MEM_DATA_IN_PRIME, ALU_OUTPUT_OUT, MEM_DATA_OUT );
  input [1:0] BYTE_LEN_IN;
  output [1:0] BYTE_LEN_OUT;
  input [31:0] ALU_OUTPUT_IN;
  input [31:0] MEM_DATA_IN;
  input [31:0] MEM_DATA_OUT_INT;
  input [31:0] NPC_IN;
  input [4:0] IR_IN;
  output [4:0] IR_OUT;
  output [31:0] NPC_OUT;
  output [31:0] MEM_ADDR_OUT;
  output [31:0] MEM_DATA_IN_PRIME;
  output [31:0] ALU_OUTPUT_OUT;
  output [31:0] MEM_DATA_OUT;
  input CLK, RST, MEM_OUTREG_EN, DRAM_WE;
  output DRAM_WE_OUT;
  wire   DRAM_WE;
  assign DRAM_WE_OUT = DRAM_WE;
  assign BYTE_LEN_OUT[1] = BYTE_LEN_IN[1];
  assign BYTE_LEN_OUT[0] = BYTE_LEN_IN[0];
  assign MEM_ADDR_OUT[31] = ALU_OUTPUT_IN[31];
  assign MEM_ADDR_OUT[30] = ALU_OUTPUT_IN[30];
  assign MEM_ADDR_OUT[29] = ALU_OUTPUT_IN[29];
  assign MEM_ADDR_OUT[28] = ALU_OUTPUT_IN[28];
  assign MEM_ADDR_OUT[27] = ALU_OUTPUT_IN[27];
  assign MEM_ADDR_OUT[26] = ALU_OUTPUT_IN[26];
  assign MEM_ADDR_OUT[25] = ALU_OUTPUT_IN[25];
  assign MEM_ADDR_OUT[24] = ALU_OUTPUT_IN[24];
  assign MEM_ADDR_OUT[23] = ALU_OUTPUT_IN[23];
  assign MEM_ADDR_OUT[22] = ALU_OUTPUT_IN[22];
  assign MEM_ADDR_OUT[21] = ALU_OUTPUT_IN[21];
  assign MEM_ADDR_OUT[20] = ALU_OUTPUT_IN[20];
  assign MEM_ADDR_OUT[19] = ALU_OUTPUT_IN[19];
  assign MEM_ADDR_OUT[18] = ALU_OUTPUT_IN[18];
  assign MEM_ADDR_OUT[17] = ALU_OUTPUT_IN[17];
  assign MEM_ADDR_OUT[16] = ALU_OUTPUT_IN[16];
  assign MEM_ADDR_OUT[15] = ALU_OUTPUT_IN[15];
  assign MEM_ADDR_OUT[14] = ALU_OUTPUT_IN[14];
  assign MEM_ADDR_OUT[13] = ALU_OUTPUT_IN[13];
  assign MEM_ADDR_OUT[12] = ALU_OUTPUT_IN[12];
  assign MEM_ADDR_OUT[11] = ALU_OUTPUT_IN[11];
  assign MEM_ADDR_OUT[10] = ALU_OUTPUT_IN[10];
  assign MEM_ADDR_OUT[9] = ALU_OUTPUT_IN[9];
  assign MEM_ADDR_OUT[8] = ALU_OUTPUT_IN[8];
  assign MEM_ADDR_OUT[7] = ALU_OUTPUT_IN[7];
  assign MEM_ADDR_OUT[6] = ALU_OUTPUT_IN[6];
  assign MEM_ADDR_OUT[5] = ALU_OUTPUT_IN[5];
  assign MEM_ADDR_OUT[4] = ALU_OUTPUT_IN[4];
  assign MEM_ADDR_OUT[3] = ALU_OUTPUT_IN[3];
  assign MEM_ADDR_OUT[2] = ALU_OUTPUT_IN[2];
  assign MEM_ADDR_OUT[1] = ALU_OUTPUT_IN[1];
  assign MEM_ADDR_OUT[0] = ALU_OUTPUT_IN[0];
  assign MEM_DATA_IN_PRIME[31] = MEM_DATA_IN[31];
  assign MEM_DATA_IN_PRIME[30] = MEM_DATA_IN[30];
  assign MEM_DATA_IN_PRIME[29] = MEM_DATA_IN[29];
  assign MEM_DATA_IN_PRIME[28] = MEM_DATA_IN[28];
  assign MEM_DATA_IN_PRIME[27] = MEM_DATA_IN[27];
  assign MEM_DATA_IN_PRIME[26] = MEM_DATA_IN[26];
  assign MEM_DATA_IN_PRIME[25] = MEM_DATA_IN[25];
  assign MEM_DATA_IN_PRIME[24] = MEM_DATA_IN[24];
  assign MEM_DATA_IN_PRIME[23] = MEM_DATA_IN[23];
  assign MEM_DATA_IN_PRIME[22] = MEM_DATA_IN[22];
  assign MEM_DATA_IN_PRIME[21] = MEM_DATA_IN[21];
  assign MEM_DATA_IN_PRIME[20] = MEM_DATA_IN[20];
  assign MEM_DATA_IN_PRIME[19] = MEM_DATA_IN[19];
  assign MEM_DATA_IN_PRIME[18] = MEM_DATA_IN[18];
  assign MEM_DATA_IN_PRIME[17] = MEM_DATA_IN[17];
  assign MEM_DATA_IN_PRIME[16] = MEM_DATA_IN[16];
  assign MEM_DATA_IN_PRIME[15] = MEM_DATA_IN[15];
  assign MEM_DATA_IN_PRIME[14] = MEM_DATA_IN[14];
  assign MEM_DATA_IN_PRIME[13] = MEM_DATA_IN[13];
  assign MEM_DATA_IN_PRIME[12] = MEM_DATA_IN[12];
  assign MEM_DATA_IN_PRIME[11] = MEM_DATA_IN[11];
  assign MEM_DATA_IN_PRIME[10] = MEM_DATA_IN[10];
  assign MEM_DATA_IN_PRIME[9] = MEM_DATA_IN[9];
  assign MEM_DATA_IN_PRIME[8] = MEM_DATA_IN[8];
  assign MEM_DATA_IN_PRIME[7] = MEM_DATA_IN[7];
  assign MEM_DATA_IN_PRIME[6] = MEM_DATA_IN[6];
  assign MEM_DATA_IN_PRIME[5] = MEM_DATA_IN[5];
  assign MEM_DATA_IN_PRIME[4] = MEM_DATA_IN[4];
  assign MEM_DATA_IN_PRIME[3] = MEM_DATA_IN[3];
  assign MEM_DATA_IN_PRIME[2] = MEM_DATA_IN[2];
  assign MEM_DATA_IN_PRIME[1] = MEM_DATA_IN[1];
  assign MEM_DATA_IN_PRIME[0] = MEM_DATA_IN[0];
  assign MEM_DATA_OUT[31] = MEM_DATA_OUT_INT[31];
  assign MEM_DATA_OUT[30] = MEM_DATA_OUT_INT[30];
  assign MEM_DATA_OUT[29] = MEM_DATA_OUT_INT[29];
  assign MEM_DATA_OUT[28] = MEM_DATA_OUT_INT[28];
  assign MEM_DATA_OUT[27] = MEM_DATA_OUT_INT[27];
  assign MEM_DATA_OUT[26] = MEM_DATA_OUT_INT[26];
  assign MEM_DATA_OUT[25] = MEM_DATA_OUT_INT[25];
  assign MEM_DATA_OUT[24] = MEM_DATA_OUT_INT[24];
  assign MEM_DATA_OUT[23] = MEM_DATA_OUT_INT[23];
  assign MEM_DATA_OUT[22] = MEM_DATA_OUT_INT[22];
  assign MEM_DATA_OUT[21] = MEM_DATA_OUT_INT[21];
  assign MEM_DATA_OUT[20] = MEM_DATA_OUT_INT[20];
  assign MEM_DATA_OUT[19] = MEM_DATA_OUT_INT[19];
  assign MEM_DATA_OUT[18] = MEM_DATA_OUT_INT[18];
  assign MEM_DATA_OUT[17] = MEM_DATA_OUT_INT[17];
  assign MEM_DATA_OUT[16] = MEM_DATA_OUT_INT[16];
  assign MEM_DATA_OUT[15] = MEM_DATA_OUT_INT[15];
  assign MEM_DATA_OUT[14] = MEM_DATA_OUT_INT[14];
  assign MEM_DATA_OUT[13] = MEM_DATA_OUT_INT[13];
  assign MEM_DATA_OUT[12] = MEM_DATA_OUT_INT[12];
  assign MEM_DATA_OUT[11] = MEM_DATA_OUT_INT[11];
  assign MEM_DATA_OUT[10] = MEM_DATA_OUT_INT[10];
  assign MEM_DATA_OUT[9] = MEM_DATA_OUT_INT[9];
  assign MEM_DATA_OUT[8] = MEM_DATA_OUT_INT[8];
  assign MEM_DATA_OUT[7] = MEM_DATA_OUT_INT[7];
  assign MEM_DATA_OUT[6] = MEM_DATA_OUT_INT[6];
  assign MEM_DATA_OUT[5] = MEM_DATA_OUT_INT[5];
  assign MEM_DATA_OUT[4] = MEM_DATA_OUT_INT[4];
  assign MEM_DATA_OUT[3] = MEM_DATA_OUT_INT[3];
  assign MEM_DATA_OUT[2] = MEM_DATA_OUT_INT[2];
  assign MEM_DATA_OUT[1] = MEM_DATA_OUT_INT[1];
  assign MEM_DATA_OUT[0] = MEM_DATA_OUT_INT[0];

  gen_reg_N32_2 PAD_ALU ( .clk(CLK), .rst(RST), .ld(MEM_OUTREG_EN), .data_in(
        ALU_OUTPUT_IN), .data_out(ALU_OUTPUT_OUT) );
  gen_reg_N32_1 NPC3 ( .clk(CLK), .rst(RST), .ld(MEM_OUTREG_EN), .data_in(
        NPC_IN), .data_out(NPC_OUT) );
  gen_reg_N5_1 IR3 ( .clk(CLK), .rst(RST), .ld(MEM_OUTREG_EN), .data_in(IR_IN), 
        .data_out(IR_OUT) );
endmodule


module gen_mux41_N32 ( sel, w, x, y, z, m );
  input [1:0] sel;
  input [31:0] w;
  input [31:0] x;
  input [31:0] y;
  input [31:0] z;
  output [31:0] m;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n74, n76, n80,
         n83, n84, n85;

  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(m[9]) );
  AOI22_X1 U4 ( .A1(w[9]), .A2(n83), .B1(x[9]), .B2(n80), .ZN(n4) );
  AOI22_X1 U5 ( .A1(y[9]), .A2(n7), .B1(z[9]), .B2(n74), .ZN(n3) );
  NAND2_X1 U6 ( .A1(n9), .A2(n10), .ZN(m[8]) );
  AOI22_X1 U7 ( .A1(w[8]), .A2(n83), .B1(x[8]), .B2(n80), .ZN(n10) );
  AOI22_X1 U8 ( .A1(y[8]), .A2(n7), .B1(z[8]), .B2(n74), .ZN(n9) );
  NAND2_X1 U9 ( .A1(n11), .A2(n12), .ZN(m[7]) );
  AOI22_X1 U10 ( .A1(w[7]), .A2(n83), .B1(x[7]), .B2(n80), .ZN(n12) );
  AOI22_X1 U11 ( .A1(y[7]), .A2(n7), .B1(z[7]), .B2(n74), .ZN(n11) );
  NAND2_X1 U12 ( .A1(n13), .A2(n14), .ZN(m[6]) );
  AOI22_X1 U13 ( .A1(w[6]), .A2(n83), .B1(x[6]), .B2(n80), .ZN(n14) );
  AOI22_X1 U14 ( .A1(y[6]), .A2(n76), .B1(z[6]), .B2(n74), .ZN(n13) );
  NAND2_X1 U15 ( .A1(n15), .A2(n16), .ZN(m[5]) );
  AOI22_X1 U16 ( .A1(w[5]), .A2(n83), .B1(x[5]), .B2(n80), .ZN(n16) );
  AOI22_X1 U17 ( .A1(y[5]), .A2(n7), .B1(z[5]), .B2(n74), .ZN(n15) );
  NAND2_X1 U18 ( .A1(n17), .A2(n18), .ZN(m[4]) );
  AOI22_X1 U19 ( .A1(w[4]), .A2(n83), .B1(x[4]), .B2(n80), .ZN(n18) );
  AOI22_X1 U20 ( .A1(y[4]), .A2(n7), .B1(z[4]), .B2(n74), .ZN(n17) );
  NAND2_X1 U21 ( .A1(n19), .A2(n20), .ZN(m[3]) );
  AOI22_X1 U22 ( .A1(w[3]), .A2(n83), .B1(x[3]), .B2(n80), .ZN(n20) );
  AOI22_X1 U23 ( .A1(y[3]), .A2(n7), .B1(z[3]), .B2(n74), .ZN(n19) );
  NAND2_X1 U24 ( .A1(n21), .A2(n22), .ZN(m[31]) );
  AOI22_X1 U25 ( .A1(w[31]), .A2(n83), .B1(x[31]), .B2(n80), .ZN(n22) );
  AOI22_X1 U26 ( .A1(y[31]), .A2(n7), .B1(z[31]), .B2(n74), .ZN(n21) );
  NAND2_X1 U27 ( .A1(n23), .A2(n24), .ZN(m[30]) );
  AOI22_X1 U28 ( .A1(w[30]), .A2(n83), .B1(x[30]), .B2(n80), .ZN(n24) );
  AOI22_X1 U29 ( .A1(y[30]), .A2(n76), .B1(z[30]), .B2(n74), .ZN(n23) );
  NAND2_X1 U30 ( .A1(n25), .A2(n26), .ZN(m[2]) );
  AOI22_X1 U31 ( .A1(w[2]), .A2(n83), .B1(x[2]), .B2(n80), .ZN(n26) );
  AOI22_X1 U32 ( .A1(y[2]), .A2(n7), .B1(z[2]), .B2(n74), .ZN(n25) );
  NAND2_X1 U33 ( .A1(n27), .A2(n28), .ZN(m[29]) );
  AOI22_X1 U34 ( .A1(w[29]), .A2(n83), .B1(x[29]), .B2(n80), .ZN(n28) );
  AOI22_X1 U35 ( .A1(y[29]), .A2(n76), .B1(z[29]), .B2(n74), .ZN(n27) );
  NAND2_X1 U36 ( .A1(n29), .A2(n30), .ZN(m[28]) );
  AOI22_X1 U37 ( .A1(w[28]), .A2(n83), .B1(x[28]), .B2(n80), .ZN(n30) );
  AOI22_X1 U38 ( .A1(y[28]), .A2(n76), .B1(z[28]), .B2(n74), .ZN(n29) );
  NAND2_X1 U39 ( .A1(n31), .A2(n32), .ZN(m[27]) );
  AOI22_X1 U40 ( .A1(w[27]), .A2(n83), .B1(x[27]), .B2(n80), .ZN(n32) );
  AOI22_X1 U41 ( .A1(y[27]), .A2(n76), .B1(z[27]), .B2(n74), .ZN(n31) );
  NAND2_X1 U42 ( .A1(n33), .A2(n34), .ZN(m[26]) );
  AOI22_X1 U43 ( .A1(w[26]), .A2(n83), .B1(x[26]), .B2(n80), .ZN(n34) );
  AOI22_X1 U44 ( .A1(y[26]), .A2(n76), .B1(z[26]), .B2(n74), .ZN(n33) );
  NAND2_X1 U45 ( .A1(n35), .A2(n36), .ZN(m[25]) );
  AOI22_X1 U46 ( .A1(w[25]), .A2(n83), .B1(x[25]), .B2(n80), .ZN(n36) );
  AOI22_X1 U47 ( .A1(y[25]), .A2(n76), .B1(z[25]), .B2(n74), .ZN(n35) );
  NAND2_X1 U48 ( .A1(n37), .A2(n38), .ZN(m[24]) );
  AOI22_X1 U49 ( .A1(w[24]), .A2(n83), .B1(x[24]), .B2(n80), .ZN(n38) );
  AOI22_X1 U50 ( .A1(y[24]), .A2(n76), .B1(z[24]), .B2(n74), .ZN(n37) );
  NAND2_X1 U51 ( .A1(n39), .A2(n40), .ZN(m[23]) );
  AOI22_X1 U52 ( .A1(w[23]), .A2(n83), .B1(x[23]), .B2(n80), .ZN(n40) );
  AOI22_X1 U53 ( .A1(y[23]), .A2(n76), .B1(z[23]), .B2(n74), .ZN(n39) );
  NAND2_X1 U54 ( .A1(n41), .A2(n42), .ZN(m[22]) );
  AOI22_X1 U55 ( .A1(w[22]), .A2(n83), .B1(x[22]), .B2(n80), .ZN(n42) );
  AOI22_X1 U56 ( .A1(y[22]), .A2(n76), .B1(z[22]), .B2(n74), .ZN(n41) );
  NAND2_X1 U57 ( .A1(n43), .A2(n44), .ZN(m[21]) );
  AOI22_X1 U58 ( .A1(w[21]), .A2(n83), .B1(x[21]), .B2(n80), .ZN(n44) );
  AOI22_X1 U59 ( .A1(y[21]), .A2(n76), .B1(z[21]), .B2(n74), .ZN(n43) );
  NAND2_X1 U60 ( .A1(n45), .A2(n46), .ZN(m[20]) );
  AOI22_X1 U61 ( .A1(w[20]), .A2(n5), .B1(x[20]), .B2(n80), .ZN(n46) );
  AOI22_X1 U62 ( .A1(y[20]), .A2(n76), .B1(z[20]), .B2(n74), .ZN(n45) );
  NAND2_X1 U63 ( .A1(n47), .A2(n48), .ZN(m[1]) );
  AOI22_X1 U64 ( .A1(w[1]), .A2(n83), .B1(x[1]), .B2(n80), .ZN(n48) );
  AOI22_X1 U65 ( .A1(y[1]), .A2(n76), .B1(z[1]), .B2(n74), .ZN(n47) );
  NAND2_X1 U66 ( .A1(n49), .A2(n50), .ZN(m[19]) );
  AOI22_X1 U67 ( .A1(w[19]), .A2(n5), .B1(x[19]), .B2(n6), .ZN(n50) );
  AOI22_X1 U68 ( .A1(y[19]), .A2(n76), .B1(z[19]), .B2(n8), .ZN(n49) );
  NAND2_X1 U69 ( .A1(n51), .A2(n52), .ZN(m[18]) );
  AOI22_X1 U70 ( .A1(w[18]), .A2(n5), .B1(x[18]), .B2(n6), .ZN(n52) );
  AOI22_X1 U71 ( .A1(y[18]), .A2(n76), .B1(z[18]), .B2(n8), .ZN(n51) );
  NAND2_X1 U72 ( .A1(n53), .A2(n54), .ZN(m[17]) );
  AOI22_X1 U73 ( .A1(w[17]), .A2(n5), .B1(x[17]), .B2(n6), .ZN(n54) );
  AOI22_X1 U74 ( .A1(y[17]), .A2(n7), .B1(z[17]), .B2(n8), .ZN(n53) );
  NAND2_X1 U75 ( .A1(n55), .A2(n56), .ZN(m[16]) );
  AOI22_X1 U76 ( .A1(w[16]), .A2(n5), .B1(x[16]), .B2(n6), .ZN(n56) );
  AOI22_X1 U77 ( .A1(y[16]), .A2(n76), .B1(z[16]), .B2(n8), .ZN(n55) );
  NAND2_X1 U78 ( .A1(n57), .A2(n58), .ZN(m[15]) );
  AOI22_X1 U79 ( .A1(w[15]), .A2(n5), .B1(x[15]), .B2(n6), .ZN(n58) );
  AOI22_X1 U80 ( .A1(y[15]), .A2(n76), .B1(z[15]), .B2(n8), .ZN(n57) );
  NAND2_X1 U81 ( .A1(n59), .A2(n60), .ZN(m[14]) );
  AOI22_X1 U82 ( .A1(w[14]), .A2(n5), .B1(x[14]), .B2(n6), .ZN(n60) );
  AOI22_X1 U83 ( .A1(y[14]), .A2(n76), .B1(z[14]), .B2(n8), .ZN(n59) );
  NAND2_X1 U84 ( .A1(n61), .A2(n62), .ZN(m[13]) );
  AOI22_X1 U85 ( .A1(w[13]), .A2(n5), .B1(x[13]), .B2(n6), .ZN(n62) );
  AOI22_X1 U86 ( .A1(y[13]), .A2(n76), .B1(z[13]), .B2(n8), .ZN(n61) );
  NAND2_X1 U87 ( .A1(n63), .A2(n64), .ZN(m[12]) );
  AOI22_X1 U88 ( .A1(w[12]), .A2(n5), .B1(x[12]), .B2(n6), .ZN(n64) );
  AOI22_X1 U89 ( .A1(y[12]), .A2(n76), .B1(z[12]), .B2(n8), .ZN(n63) );
  NAND2_X1 U90 ( .A1(n65), .A2(n66), .ZN(m[11]) );
  AOI22_X1 U91 ( .A1(w[11]), .A2(n5), .B1(x[11]), .B2(n6), .ZN(n66) );
  AOI22_X1 U92 ( .A1(y[11]), .A2(n76), .B1(z[11]), .B2(n8), .ZN(n65) );
  NAND2_X1 U93 ( .A1(n67), .A2(n68), .ZN(m[10]) );
  AOI22_X1 U94 ( .A1(w[10]), .A2(n83), .B1(x[10]), .B2(n80), .ZN(n68) );
  AOI22_X1 U95 ( .A1(y[10]), .A2(n76), .B1(z[10]), .B2(n8), .ZN(n67) );
  NAND2_X1 U96 ( .A1(n69), .A2(n70), .ZN(m[0]) );
  AOI22_X1 U97 ( .A1(w[0]), .A2(n83), .B1(x[0]), .B2(n6), .ZN(n70) );
  NOR2_X1 U98 ( .A1(n85), .A2(sel[1]), .ZN(n6) );
  NOR2_X1 U99 ( .A1(sel[0]), .A2(sel[1]), .ZN(n5) );
  AOI22_X1 U100 ( .A1(y[0]), .A2(n7), .B1(z[0]), .B2(n74), .ZN(n69) );
  NOR2_X1 U101 ( .A1(n84), .A2(n85), .ZN(n8) );
  NOR2_X1 U102 ( .A1(n84), .A2(sel[0]), .ZN(n7) );
  CLKBUF_X1 U103 ( .A(n8), .Z(n74) );
  CLKBUF_X1 U106 ( .A(n7), .Z(n76) );
  CLKBUF_X1 U111 ( .A(n5), .Z(n83) );
  CLKBUF_X1 U112 ( .A(n6), .Z(n80) );
  INV_X1 U113 ( .A(sel[1]), .ZN(n84) );
  INV_X1 U114 ( .A(sel[0]), .ZN(n85) );
endmodule


module sign_ext_alt_N_IN016_N_IN18_N_OUT32 ( ctrl_in, zero_padding, data_in, 
        data_ext );
  input [15:0] data_in;
  output [31:0] data_ext;
  input ctrl_in, zero_padding;
  wire   \data_ext[31] , \data_in[7] , \data_in[6] , \data_in[5] ,
         \data_in[4] , \data_in[3] , \data_in[2] , \data_in[1] , \data_in[0] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, \data_ext[30] , n16, n17;
  assign data_ext[23] = \data_ext[31] ;
  assign data_ext[17] = \data_ext[31] ;
  assign data_ext[16] = \data_ext[31] ;
  assign data_ext[22] = \data_ext[31] ;
  assign data_ext[25] = \data_ext[31] ;
  assign data_ext[31] = \data_ext[31] ;
  assign data_ext[7] = \data_in[7] ;
  assign \data_in[7]  = data_in[7];
  assign data_ext[6] = \data_in[6] ;
  assign \data_in[6]  = data_in[6];
  assign data_ext[5] = \data_in[5] ;
  assign \data_in[5]  = data_in[5];
  assign data_ext[4] = \data_in[4] ;
  assign \data_in[4]  = data_in[4];
  assign data_ext[3] = \data_in[3] ;
  assign \data_in[3]  = data_in[3];
  assign data_ext[2] = \data_in[2] ;
  assign \data_in[2]  = data_in[2];
  assign data_ext[1] = \data_in[1] ;
  assign \data_in[1]  = data_in[1];
  assign data_ext[0] = \data_in[0] ;
  assign \data_in[0]  = data_in[0];
  assign data_ext[29] = \data_ext[30] ;
  assign data_ext[26] = \data_ext[30] ;
  assign data_ext[20] = \data_ext[30] ;
  assign data_ext[19] = \data_ext[30] ;
  assign data_ext[28] = \data_ext[30] ;
  assign data_ext[18] = \data_ext[30] ;
  assign data_ext[21] = \data_ext[30] ;
  assign data_ext[24] = \data_ext[30] ;
  assign data_ext[27] = \data_ext[30] ;
  assign data_ext[30] = \data_ext[30] ;

  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(data_ext[9]) );
  NAND2_X1 U5 ( .A1(data_in[9]), .A2(ctrl_in), .ZN(n4) );
  NAND2_X1 U6 ( .A1(n3), .A2(n5), .ZN(data_ext[8]) );
  NAND2_X1 U7 ( .A1(data_in[8]), .A2(ctrl_in), .ZN(n5) );
  OAI21_X1 U8 ( .B1(n17), .B2(n6), .A(n3), .ZN(\data_ext[31] ) );
  OR2_X1 U9 ( .A1(n16), .A2(zero_padding), .ZN(n6) );
  OAI21_X1 U10 ( .B1(n16), .B2(n17), .A(n3), .ZN(data_ext[15]) );
  NAND2_X1 U11 ( .A1(n3), .A2(n7), .ZN(data_ext[14]) );
  NAND2_X1 U12 ( .A1(data_in[14]), .A2(ctrl_in), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n3), .A2(n8), .ZN(data_ext[13]) );
  NAND2_X1 U14 ( .A1(data_in[13]), .A2(ctrl_in), .ZN(n8) );
  NAND2_X1 U15 ( .A1(n3), .A2(n9), .ZN(data_ext[12]) );
  NAND2_X1 U16 ( .A1(data_in[12]), .A2(ctrl_in), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n3), .A2(n10), .ZN(data_ext[11]) );
  NAND2_X1 U18 ( .A1(data_in[11]), .A2(ctrl_in), .ZN(n10) );
  NAND2_X1 U19 ( .A1(n3), .A2(n11), .ZN(data_ext[10]) );
  NAND2_X1 U20 ( .A1(data_in[10]), .A2(ctrl_in), .ZN(n11) );
  NAND2_X1 U21 ( .A1(n12), .A2(\data_in[7] ), .ZN(n3) );
  NOR2_X1 U22 ( .A1(zero_padding), .A2(ctrl_in), .ZN(n12) );
  CLKBUF_X1 U23 ( .A(\data_ext[31] ), .Z(\data_ext[30] ) );
  INV_X1 U24 ( .A(ctrl_in), .ZN(n16) );
  INV_X1 U25 ( .A(data_in[15]), .ZN(n17) );
endmodule


module WB_STAGE_N_BITS_DATA32 ( WB_MUX_SEL, WB_CTRL_SIGN, ZERO_PADDING5, 
        NPC_OUT, MEM_OUT, ALU_OUT, MUX_OUT );
  input [1:0] WB_MUX_SEL;
  input [31:0] NPC_OUT;
  input [31:0] MEM_OUT;
  input [31:0] ALU_OUT;
  output [31:0] MUX_OUT;
  input WB_CTRL_SIGN, ZERO_PADDING5;

  wire   [31:0] SIGN_OUT;

  gen_mux41_N32 MUX ( .sel(WB_MUX_SEL), .w(ALU_OUT), .x(MEM_OUT), .y(SIGN_OUT), 
        .z(NPC_OUT), .m(MUX_OUT) );
  sign_ext_alt_N_IN016_N_IN18_N_OUT32 SIGN_EXTEND ( .ctrl_in(WB_CTRL_SIGN), 
        .zero_padding(ZERO_PADDING5), .data_in(MEM_OUT[15:0]), .data_ext(
        SIGN_OUT) );
endmodule


module DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 ( 
        CLK, RST, IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, WR_EN, 
        JAL_REG31, ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, 
        JUMP_EN, .ALU_OPCODE({\ALU_OPCODE[6] , \ALU_OPCODE[5] , 
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), MEM_OUTREG_EN, BYTE_LEN_IN, DRAM_WE, DRAM_WE_OUT, 
        BYTE_LEN_OUT, WB_MUX_SEL, WB_CTRL_SIGN, ZERO_PADDING5, IR_IN, PC_OUT, 
        MEM_DATA_OUT_INT, MEM_ADDR_OUT, MEM_DATA_IN_PRIME );
  input [1:0] BYTE_LEN_IN;
  output [1:0] BYTE_LEN_OUT;
  input [1:0] WB_MUX_SEL;
  input [31:0] IR_IN;
  output [31:0] PC_OUT;
  input [31:0] MEM_DATA_OUT_INT;
  output [31:0] MEM_ADDR_OUT;
  output [31:0] MEM_DATA_IN_PRIME;
  input CLK, RST, IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, WR_EN,
         JAL_REG31, ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND,
         JUMP_EN, \ALU_OPCODE[6] , \ALU_OPCODE[5] , \ALU_OPCODE[4] ,
         \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] ,
         MEM_OUTREG_EN, DRAM_WE, WB_CTRL_SIGN, ZERO_PADDING5;
  output DRAM_WE_OUT;

  wire   [6:0] ALU_OPCODE;
  wire   [31:0] PC_EXE2IF;
  wire   [31:0] IR_IF2ID;
  wire   [31:0] NPC_IF2EXE;
  wire   [31:0] NPC_IF2ID;
  wire   [31:0] MUX_WB2ID;
  wire   [4:0] IR_MEM2ID;
  wire   [31:0] A_ID2EXE;
  wire   [31:0] B_ID2EXE;
  wire   [31:0] IMM_ID2EXE;
  wire   [4:0] IR_ID2EXE;
  wire   [31:0] NPC_ID2EXE;
  wire   [31:0] NPC_EXE2MEM;
  wire   [31:0] ALU_EXE2MEM;
  wire   [31:0] PAD_EXE2MEM;
  wire   [4:0] IR_EXE2MEM;
  wire   [31:0] NPC_MEM2WB;
  wire   [31:0] ALU_MEM2WB;
  wire   [31:0] MEM_MEM2WB;

  IF_STAGE_N_BITS_DATA32_N_BYTES_INST4 FETCH ( .CLK(CLK), .RST(RST), 
        .IF_LATCH_EN(IF_LATCH_EN), .PC_IN(PC_EXE2IF), .IR_IN(IR_IN), .PC_OUT(
        PC_OUT), .IR_OUT(IR_IF2ID), .ADD_OUT(NPC_IF2EXE), .NPC_OUT(NPC_IF2ID)
         );
  ID_STAGE_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 DECODE ( 
        .CLK(CLK), .RST(RST), .JAL_REG31(JAL_REG31), .DEC_OUTREG_EN(
        DEC_OUTREG_EN), .IS_I_TYPE(IS_I_TYPE), .RD1_EN(RD1_EN), .RD2_EN(RD2_EN), .WR_EN(WR_EN), .ZERO_PADDING2(ZERO_PADDING2), .I_CODE(IR_IF2ID), .NPC1_IN(
        NPC_IF2ID), .DATA_IN(MUX_WB2ID), .WR_ADDR_IN(IR_MEM2ID), .REGA_OUT(
        A_ID2EXE), .REGB_OUT(B_ID2EXE), .REGIMM_OUT(IMM_ID2EXE), .WR_ADDR_OUT(
        IR_ID2EXE), .NPC1_OUT(NPC_ID2EXE) );
  EXE_STAGE_N_BITS_DATA32_RF_ADDR5 EXECUTE ( .CLK(CLK), .RST(RST), .MUXA_SEL(
        MUXA_SEL), .MUXB_SEL(MUXB_SEL), .EXE_OUTREG_EN(EXE_OUTREG_EN), 
        .EQ_COND(EQ_COND), .JUMP_EN(JUMP_EN), .ALU_OPCODE({\ALU_OPCODE[6] , 
        \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , 
        \ALU_OPCODE[1] , \ALU_OPCODE[0] }), .NPC2_IN(NPC_ID2EXE), 
        .NPC1_MUXA_IN(NPC_ID2EXE), .REGA_MUXA_IN(A_ID2EXE), .REGB_MUXB_IN(
        B_ID2EXE), .IMM_MUXB_IN(IMM_ID2EXE), .PAD_IN(B_ID2EXE), .IR2_IN(
        IR_ID2EXE), .JUMP_MUX_IN_0(NPC_IF2EXE), .NPC2_OUT(NPC_EXE2MEM), 
        .ALU_OUT(ALU_EXE2MEM), .PAD_OUT(PAD_EXE2MEM), .IR2_OUT(IR_EXE2MEM), 
        .ADDR_MUX_OUT(PC_EXE2IF) );
  MEM_STAGE_N_BITS_DATA32_RF_ADDR5 MEMORY ( .CLK(CLK), .RST(RST), 
        .MEM_OUTREG_EN(MEM_OUTREG_EN), .BYTE_LEN_IN(BYTE_LEN_IN), .DRAM_WE(
        DRAM_WE), .DRAM_WE_OUT(DRAM_WE_OUT), .BYTE_LEN_OUT(BYTE_LEN_OUT), 
        .ALU_OUTPUT_IN(ALU_EXE2MEM), .MEM_DATA_IN(PAD_EXE2MEM), 
        .MEM_DATA_OUT_INT(MEM_DATA_OUT_INT), .NPC_IN(NPC_EXE2MEM), .IR_IN(
        IR_EXE2MEM), .IR_OUT(IR_MEM2ID), .NPC_OUT(NPC_MEM2WB), .MEM_ADDR_OUT(
        MEM_ADDR_OUT), .MEM_DATA_IN_PRIME(MEM_DATA_IN_PRIME), .ALU_OUTPUT_OUT(
        ALU_MEM2WB), .MEM_DATA_OUT(MEM_MEM2WB) );
  WB_STAGE_N_BITS_DATA32 WRITE_BACK ( .WB_MUX_SEL(WB_MUX_SEL), .WB_CTRL_SIGN(
        WB_CTRL_SIGN), .ZERO_PADDING5(ZERO_PADDING5), .NPC_OUT(NPC_MEM2WB), 
        .MEM_OUT(MEM_MEM2WB), .ALU_OUT(ALU_MEM2WB), .MUX_OUT(MUX_WB2ID) );
endmodule


module CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE20 ( Clk, 
        Rst, IR_IN, IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, 
        ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN, 
    .ALU_OPCODE({\ALU_OPCODE[6] , \ALU_OPCODE[5] , \ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), 
    .FPU_OPCODE({\FPU_OPCODE[4] , \FPU_OPCODE[3] , \FPU_OPCODE[2] , 
        \FPU_OPCODE[1] , \FPU_OPCODE[0] }), MEM_OUTREG_EN, DRAM_WE, BYTE_LEN, 
        WB_MUX_SEL, JAL_REG31, WB_CTRL_SIGN, ZERO_PADDING5, WR_EN );
  input [31:0] IR_IN;
  output [1:0] BYTE_LEN;
  output [1:0] WB_MUX_SEL;
  input Clk, Rst;
  output IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, ZERO_PADDING2,
         MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND, JUMP_EN, \ALU_OPCODE[6] ,
         \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] ,
         \ALU_OPCODE[1] , \ALU_OPCODE[0] , \FPU_OPCODE[4] , \FPU_OPCODE[3] ,
         \FPU_OPCODE[2] , \FPU_OPCODE[1] , \FPU_OPCODE[0] , MEM_OUTREG_EN,
         DRAM_WE, JAL_REG31, WB_CTRL_SIGN, ZERO_PADDING5, WR_EN;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26,
         \ALU_op[5] , n26, n38, n46, n57, n63, n82, n315, n327, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n243, n244, n245, n246, n247, n248, n249,
         n252, n253, n254, n275, n276, n277, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n317, n318,
         n319, n320, n322, n323, n324, n325, n326, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337;
  wire   [6:0] ALU_OPCODE;
  wire   [4:0] FPU_OPCODE;
  wire   [18:0] cw1;
  wire   [13:0] cw2;
  wire   [8:0] cw3;
  wire   [4:0] cw4;
  wire   [6:0] ALU_op1;
  wire   [6:0] ALU_op2;
  wire   [4:0] FPU_op1;
  wire   [4:0] FPU_op2;
  wire   [19:0] cw;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];

  OAI21_X1 U67 ( .B1(n276), .B2(n64), .A(n65), .ZN(n252) );
  NOR2_X1 U68 ( .A1(n66), .A2(n293), .ZN(n65) );
  NAND2_X1 U69 ( .A1(n68), .A2(n69), .ZN(n82) );
  AOI21_X1 U70 ( .B1(n70), .B2(n71), .A(n72), .ZN(n69) );
  AOI21_X1 U71 ( .B1(n296), .B2(IR_IN_31), .A(n307), .ZN(n72) );
  AOI21_X1 U72 ( .B1(n74), .B2(n75), .A(IR_IN_28), .ZN(n70) );
  NOR4_X1 U73 ( .A1(n76), .A2(n318), .A3(n77), .A4(n78), .ZN(n75) );
  NOR2_X1 U74 ( .A1(n79), .A2(n311), .ZN(n78) );
  AOI21_X1 U75 ( .B1(n80), .B2(n325), .A(n317), .ZN(n77) );
  AOI21_X1 U77 ( .B1(n84), .B2(n85), .A(n86), .ZN(n83) );
  AOI22_X1 U78 ( .A1(IR_IN_31), .A2(n87), .B1(n303), .B2(n295), .ZN(n68) );
  OAI21_X1 U79 ( .B1(IR_IN_27), .B2(n88), .A(n89), .ZN(n87) );
  AOI22_X1 U80 ( .A1(n295), .A2(n90), .B1(n91), .B2(n92), .ZN(n88) );
  OR2_X1 U81 ( .A1(n93), .A2(n94), .ZN(n63) );
  OAI21_X1 U82 ( .B1(n95), .B2(n304), .A(n96), .ZN(n94) );
  AOI22_X1 U83 ( .A1(n289), .A2(n97), .B1(n303), .B2(n71), .ZN(n96) );
  OAI21_X1 U84 ( .B1(n99), .B2(n100), .A(n101), .ZN(n93) );
  AOI21_X1 U85 ( .B1(n102), .B2(n335), .A(n287), .ZN(n101) );
  OAI21_X1 U86 ( .B1(n103), .B2(n282), .A(n104), .ZN(n57) );
  AOI21_X1 U87 ( .B1(n105), .B2(n299), .A(n106), .ZN(n104) );
  NOR3_X1 U88 ( .A1(n299), .A2(n283), .A3(n304), .ZN(n106) );
  OAI21_X1 U89 ( .B1(IR_IN_28), .B2(n107), .A(n108), .ZN(n105) );
  NOR3_X1 U90 ( .A1(n109), .A2(n110), .A3(n111), .ZN(n107) );
  OAI21_X1 U91 ( .B1(n79), .B2(n314), .A(n112), .ZN(n109) );
  NOR2_X1 U92 ( .A1(IR_IN_30), .A2(n113), .ZN(n112) );
  AOI22_X1 U93 ( .A1(n114), .A2(n115), .B1(IR_IN_30), .B2(n90), .ZN(n103) );
  NAND2_X1 U94 ( .A1(n305), .A2(IR_IN_26), .ZN(n115) );
  OAI21_X1 U95 ( .B1(n90), .B2(n116), .A(IR_IN_29), .ZN(n114) );
  NAND2_X1 U96 ( .A1(IR_IN_27), .A2(n297), .ZN(n116) );
  NOR3_X1 U98 ( .A1(n100), .A2(n307), .A3(n99), .ZN(n120) );
  OAI33_X1 U99 ( .A1(n294), .A2(IR_IN_31), .A3(IR_IN_28), .B1(n92), .B2(n282), 
        .B3(n97), .ZN(n119) );
  OAI21_X1 U100 ( .B1(n254), .B2(n304), .A(n121), .ZN(n118) );
  AOI22_X1 U101 ( .A1(n102), .A2(n122), .B1(n285), .B2(n300), .ZN(n121) );
  NAND2_X1 U102 ( .A1(n312), .A2(n123), .ZN(n122) );
  NAND2_X1 U103 ( .A1(n125), .A2(n126), .ZN(n46) );
  AOI21_X1 U104 ( .B1(n127), .B2(n282), .A(n128), .ZN(n126) );
  NOR3_X1 U105 ( .A1(n98), .A2(n300), .A3(n307), .ZN(n128) );
  OR2_X1 U106 ( .A1(n129), .A2(IR_IN_26), .ZN(n127) );
  NOR4_X1 U107 ( .A1(IR_IN_28), .A2(IR_IN_27), .A3(n130), .A4(n131), .ZN(n129)
         );
  NOR3_X1 U108 ( .A1(n132), .A2(n110), .A3(n133), .ZN(n130) );
  OAI21_X1 U109 ( .B1(n79), .B2(n317), .A(n134), .ZN(n133) );
  OAI21_X1 U110 ( .B1(n135), .B2(n81), .A(n84), .ZN(n134) );
  NAND2_X1 U111 ( .A1(n136), .A2(n137), .ZN(n110) );
  NOR3_X1 U112 ( .A1(n310), .A2(n138), .A3(n145), .ZN(n137) );
  OAI21_X1 U113 ( .B1(n326), .B2(n85), .A(n111), .ZN(n146) );
  NAND2_X1 U114 ( .A1(n311), .A2(n147), .ZN(n111) );
  AOI21_X1 U115 ( .B1(n330), .B2(n84), .A(n148), .ZN(n136) );
  OAI21_X1 U116 ( .B1(n323), .B2(n320), .A(n149), .ZN(n132) );
  NOR2_X1 U117 ( .A1(n150), .A2(n318), .ZN(n149) );
  OAI21_X1 U118 ( .B1(n152), .B2(n85), .A(n153), .ZN(n151) );
  AOI22_X1 U119 ( .A1(n283), .A2(n73), .B1(IR_IN_31), .B2(n154), .ZN(n125) );
  OAI21_X1 U120 ( .B1(IR_IN_27), .B2(n155), .A(n156), .ZN(n154) );
  AOI21_X1 U121 ( .B1(n157), .B2(n295), .A(n298), .ZN(n156) );
  NOR2_X1 U122 ( .A1(n306), .A2(n307), .ZN(n157) );
  AOI22_X1 U123 ( .A1(n301), .A2(n92), .B1(n295), .B2(n158), .ZN(n155) );
  OAI21_X1 U124 ( .B1(n302), .B2(n297), .A(n159), .ZN(n73) );
  NAND2_X1 U125 ( .A1(n309), .A2(n299), .ZN(n159) );
  OAI21_X1 U126 ( .B1(n294), .B2(n282), .A(n160), .ZN(n38) );
  AOI22_X1 U127 ( .A1(n161), .A2(n162), .B1(n283), .B2(n100), .ZN(n160) );
  OAI21_X1 U128 ( .B1(n309), .B2(n304), .A(n90), .ZN(n100) );
  OAI21_X1 U129 ( .B1(IR_IN_28), .B2(n164), .A(n98), .ZN(n162) );
  OAI21_X1 U130 ( .B1(IR_IN_30), .B2(n308), .A(n97), .ZN(n161) );
  NAND2_X1 U131 ( .A1(n309), .A2(n165), .ZN(n148) );
  NAND2_X1 U132 ( .A1(n166), .A2(n167), .ZN(n165) );
  NOR3_X1 U133 ( .A1(n168), .A2(n169), .A3(n150), .ZN(n167) );
  NOR3_X1 U134 ( .A1(n170), .A2(IR_IN[3]), .A3(n319), .ZN(n168) );
  NOR3_X1 U135 ( .A1(n86), .A2(n124), .A3(n335), .ZN(n166) );
  OAI21_X1 U137 ( .B1(n173), .B2(n147), .A(n123), .ZN(n172) );
  NOR2_X1 U138 ( .A1(n174), .A2(n175), .ZN(n123) );
  AOI21_X1 U139 ( .B1(n176), .B2(n177), .A(n317), .ZN(n175) );
  NOR2_X1 U140 ( .A1(n178), .A2(n179), .ZN(n153) );
  NAND2_X1 U141 ( .A1(n324), .A2(IR_IN[5]), .ZN(n178) );
  OAI21_X1 U142 ( .B1(n180), .B2(n314), .A(n181), .ZN(n124) );
  AOI22_X1 U143 ( .A1(n182), .A2(n183), .B1(n184), .B2(n185), .ZN(n181) );
  NAND2_X1 U144 ( .A1(n180), .A2(n79), .ZN(n185) );
  NOR2_X1 U145 ( .A1(IR_IN[3]), .A2(n186), .ZN(n182) );
  NOR2_X1 U147 ( .A1(n85), .A2(n81), .ZN(n173) );
  NOR2_X1 U148 ( .A1(n187), .A2(IR_IN[0]), .ZN(n81) );
  NOR2_X1 U149 ( .A1(n187), .A2(n333), .ZN(n85) );
  OAI21_X1 U150 ( .B1(n188), .B2(n332), .A(n189), .ZN(n86) );
  AOI21_X1 U151 ( .B1(n190), .B2(n152), .A(n138), .ZN(n189) );
  NOR2_X1 U152 ( .A1(n191), .A2(n320), .ZN(n138) );
  NOR4_X1 U153 ( .A1(IR_IN[2]), .A2(IR_IN[1]), .A3(n334), .A4(n333), .ZN(n183)
         );
  OR2_X1 U154 ( .A1(n186), .A2(n324), .ZN(n191) );
  NOR2_X1 U155 ( .A1(IR_IN[3]), .A2(n319), .ZN(n190) );
  OAI21_X1 U157 ( .B1(n324), .B2(n193), .A(n253), .ZN(n192) );
  NOR4_X1 U158 ( .A1(IR_IN[6]), .A2(IR_IN[5]), .A3(n334), .A4(n194), .ZN(n253)
         );
  NAND2_X1 U159 ( .A1(n290), .A2(n195), .ZN(n26) );
  AOI22_X1 U160 ( .A1(n306), .A2(n292), .B1(n303), .B2(n71), .ZN(n196) );
  OAI21_X1 U161 ( .B1(IR_IN_29), .B2(n197), .A(n198), .ZN(cw[9]) );
  NAND2_X1 U162 ( .A1(n286), .A2(n292), .ZN(n198) );
  NOR3_X1 U163 ( .A1(n163), .A2(IR_IN_30), .A3(n158), .ZN(cw[6]) );
  NAND2_X1 U164 ( .A1(IR_IN_31), .A2(IR_IN_27), .ZN(n163) );
  AOI21_X1 U165 ( .B1(IR_IN_26), .B2(n287), .A(n201), .ZN(n200) );
  NOR3_X1 U166 ( .A1(n282), .A2(IR_IN_30), .A3(n158), .ZN(n201) );
  OAI21_X1 U167 ( .B1(IR_IN_28), .B2(n254), .A(n284), .ZN(cw[4]) );
  OAI21_X1 U168 ( .B1(n254), .B2(n304), .A(n202), .ZN(cw[3]) );
  NOR2_X1 U169 ( .A1(cw[2]), .A2(n203), .ZN(n202) );
  NOR4_X1 U170 ( .A1(IR_IN_31), .A2(IR_IN_29), .A3(n307), .A4(n158), .ZN(cw[2]) );
  NAND2_X1 U171 ( .A1(n199), .A2(n204), .ZN(cw[15]) );
  NAND2_X1 U172 ( .A1(n205), .A2(n295), .ZN(n199) );
  NOR2_X1 U173 ( .A1(n206), .A2(n282), .ZN(n205) );
  NAND2_X1 U174 ( .A1(n207), .A2(n208), .ZN(cw[14]) );
  AOI22_X1 U175 ( .A1(n285), .A2(n209), .B1(n275), .B2(n210), .ZN(n208) );
  NAND2_X1 U176 ( .A1(n91), .A2(n97), .ZN(n210) );
  OAI21_X1 U177 ( .B1(IR_IN_27), .B2(n304), .A(n108), .ZN(n209) );
  AOI22_X1 U178 ( .A1(n212), .A2(n90), .B1(n169), .B2(n102), .ZN(n207) );
  NAND2_X1 U179 ( .A1(n213), .A2(n214), .ZN(cw[13]) );
  NOR2_X1 U180 ( .A1(n66), .A2(n215), .ZN(n214) );
  AOI21_X1 U181 ( .B1(n102), .B2(n216), .A(n217), .ZN(n213) );
  OAI21_X1 U182 ( .B1(n331), .B2(n188), .A(n313), .ZN(n216) );
  AOI21_X1 U183 ( .B1(n327), .B2(n219), .A(n64), .ZN(cw[12]) );
  OAI21_X1 U184 ( .B1(n211), .B2(n97), .A(n220), .ZN(n64) );
  NOR2_X1 U185 ( .A1(n102), .A2(n290), .ZN(n220) );
  NAND2_X1 U186 ( .A1(n302), .A2(n292), .ZN(n194) );
  NAND2_X1 U187 ( .A1(n221), .A2(IR_IN_31), .ZN(n211) );
  NOR2_X1 U188 ( .A1(n297), .A2(n299), .ZN(n221) );
  NAND2_X1 U189 ( .A1(n279), .A2(n297), .ZN(n219) );
  NAND2_X1 U190 ( .A1(n303), .A2(n282), .ZN(n197) );
  AOI21_X1 U191 ( .B1(IR_IN_28), .B2(n66), .A(n67), .ZN(n327) );
  NAND2_X1 U192 ( .A1(n222), .A2(n223), .ZN(n67) );
  AOI21_X1 U193 ( .B1(n224), .B2(n307), .A(n215), .ZN(n222) );
  NOR2_X1 U194 ( .A1(n225), .A2(n282), .ZN(n215) );
  OR2_X1 U195 ( .A1(IR_IN_30), .A2(n206), .ZN(n225) );
  AOI21_X1 U196 ( .B1(n304), .B2(n307), .A(n302), .ZN(n206) );
  OAI21_X1 U197 ( .B1(IR_IN_31), .B2(n91), .A(n131), .ZN(n224) );
  NAND2_X1 U199 ( .A1(n228), .A2(n223), .ZN(n217) );
  AOI21_X1 U200 ( .B1(n277), .B2(IR_IN_29), .A(n212), .ZN(n223) );
  AOI22_X1 U201 ( .A1(IR_IN_30), .A2(n230), .B1(n97), .B2(n282), .ZN(n229) );
  OAI21_X1 U202 ( .B1(n305), .B2(n304), .A(n108), .ZN(n230) );
  NAND2_X1 U203 ( .A1(IR_IN_27), .A2(n304), .ZN(n108) );
  NAND2_X1 U204 ( .A1(IR_IN_28), .A2(IR_IN_27), .ZN(n97) );
  AOI21_X1 U205 ( .B1(n306), .B2(n275), .A(n287), .ZN(n228) );
  NOR2_X1 U207 ( .A1(n307), .A2(n95), .ZN(n66) );
  OAI21_X1 U208 ( .B1(n231), .B2(n218), .A(n102), .ZN(n204) );
  NOR2_X1 U209 ( .A1(n90), .A2(n164), .ZN(n102) );
  NAND2_X1 U210 ( .A1(n71), .A2(n307), .ZN(n164) );
  NAND2_X1 U211 ( .A1(n232), .A2(n233), .ZN(n218) );
  NOR3_X1 U212 ( .A1(n150), .A2(n169), .A3(n76), .ZN(n233) );
  AOI21_X1 U213 ( .B1(n170), .B2(n79), .A(n147), .ZN(n76) );
  NOR2_X1 U214 ( .A1(n314), .A2(n177), .ZN(n169) );
  NOR2_X1 U215 ( .A1(n326), .A2(n330), .ZN(n177) );
  NAND2_X1 U216 ( .A1(n234), .A2(IR_IN[0]), .ZN(n79) );
  NOR2_X1 U217 ( .A1(IR_IN[1]), .A2(n328), .ZN(n234) );
  NOR2_X1 U218 ( .A1(n235), .A2(n319), .ZN(n150) );
  NAND2_X1 U219 ( .A1(n324), .A2(n330), .ZN(n235) );
  NOR3_X1 U220 ( .A1(n174), .A2(n236), .A3(n237), .ZN(n232) );
  NOR2_X1 U221 ( .A1(n147), .A2(n187), .ZN(n237) );
  NAND2_X1 U222 ( .A1(IR_IN[1]), .A2(n328), .ZN(n187) );
  NAND2_X1 U223 ( .A1(n238), .A2(IR_IN[3]), .ZN(n147) );
  NOR2_X1 U224 ( .A1(n322), .A2(n179), .ZN(n238) );
  NOR3_X1 U225 ( .A1(n319), .A2(IR_IN[3]), .A3(n176), .ZN(n236) );
  NOR2_X1 U226 ( .A1(n329), .A2(n152), .ZN(n176) );
  NOR2_X1 U227 ( .A1(n333), .A2(n193), .ZN(n152) );
  NAND2_X1 U228 ( .A1(n135), .A2(IR_IN[2]), .ZN(n170) );
  NOR2_X1 U229 ( .A1(IR_IN[0]), .A2(IR_IN[1]), .ZN(n135) );
  OR2_X1 U230 ( .A1(n145), .A2(n113), .ZN(n174) );
  NOR2_X1 U231 ( .A1(n239), .A2(n319), .ZN(n113) );
  NOR4_X1 U232 ( .A1(IR_IN[6]), .A2(IR_IN[5]), .A3(IR_IN[4]), .A4(n334), .ZN(
        n195) );
  NAND2_X1 U233 ( .A1(IR_IN[3]), .A2(n330), .ZN(n239) );
  NOR4_X1 U234 ( .A1(IR_IN[5]), .A2(IR_IN[3]), .A3(n179), .A4(n80), .ZN(n145)
         );
  NAND2_X1 U235 ( .A1(n331), .A2(n333), .ZN(n80) );
  NAND2_X1 U236 ( .A1(n240), .A2(IR_IN[4]), .ZN(n179) );
  NOR2_X1 U237 ( .A1(IR_IN[6]), .A2(n334), .ZN(n240) );
  AOI21_X1 U238 ( .B1(n311), .B2(n314), .A(n331), .ZN(n231) );
  NAND2_X1 U239 ( .A1(IR_IN[2]), .A2(IR_IN[1]), .ZN(n193) );
  NOR2_X1 U240 ( .A1(n188), .A2(IR_IN[3]), .ZN(n84) );
  NOR2_X1 U241 ( .A1(n324), .A2(n188), .ZN(n184) );
  OR2_X1 U242 ( .A1(n334), .A2(n186), .ZN(n188) );
  NAND2_X1 U243 ( .A1(n241), .A2(IR_IN[5]), .ZN(n186) );
  NOR2_X1 U244 ( .A1(IR_IN[6]), .A2(IR_IN[4]), .ZN(n241) );
  NOR2_X1 U246 ( .A1(n243), .A2(n158), .ZN(n203) );
  NAND2_X1 U247 ( .A1(IR_IN_27), .A2(n294), .ZN(n243) );
  NAND2_X1 U248 ( .A1(n244), .A2(n245), .ZN(\ALU_op[5] ) );
  NOR3_X1 U249 ( .A1(n212), .A2(n275), .A3(n287), .ZN(n245) );
  NAND2_X1 U250 ( .A1(n288), .A2(n307), .ZN(n254) );
  NAND2_X1 U251 ( .A1(n298), .A2(n282), .ZN(n95) );
  NAND2_X1 U252 ( .A1(IR_IN_30), .A2(n299), .ZN(n89) );
  NOR2_X1 U253 ( .A1(n92), .A2(IR_IN_31), .ZN(n212) );
  NAND2_X1 U254 ( .A1(IR_IN_29), .A2(n297), .ZN(n92) );
  AOI21_X1 U255 ( .B1(IR_IN_28), .B2(n71), .A(n246), .ZN(n244) );
  OAI21_X1 U256 ( .B1(n247), .B2(n98), .A(n248), .ZN(n246) );
  OAI21_X1 U257 ( .B1(n302), .B2(n306), .A(n288), .ZN(n248) );
  NAND2_X1 U258 ( .A1(IR_IN_31), .A2(n294), .ZN(n99) );
  NAND2_X1 U259 ( .A1(IR_IN_28), .A2(n309), .ZN(n91) );
  NAND2_X1 U260 ( .A1(n249), .A2(IR_IN_29), .ZN(n98) );
  NOR2_X1 U261 ( .A1(IR_IN_31), .A2(n297), .ZN(n249) );
  NOR3_X1 U262 ( .A1(n307), .A2(n300), .A3(n302), .ZN(n247) );
  NAND2_X1 U263 ( .A1(IR_IN_26), .A2(n304), .ZN(n158) );
  NAND2_X1 U264 ( .A1(n309), .A2(n304), .ZN(n90) );
  NOR2_X1 U265 ( .A1(n131), .A2(IR_IN_31), .ZN(n71) );
  NAND2_X1 U266 ( .A1(n299), .A2(n297), .ZN(n131) );
  INV_X1 U13 ( .A(n204), .ZN(n293) );
  INV_X1 U14 ( .A(n194), .ZN(n290) );
  INV_X1 U15 ( .A(n90), .ZN(n300) );
  INV_X1 U16 ( .A(n254), .ZN(n287) );
  INV_X1 U17 ( .A(n131), .ZN(n294) );
  INV_X1 U18 ( .A(n164), .ZN(n292) );
  INV_X1 U19 ( .A(n80), .ZN(n330) );
  INV_X1 U20 ( .A(n100), .ZN(n301) );
  INV_X1 U21 ( .A(n95), .ZN(n275) );
  INV_X1 U22 ( .A(n64), .ZN(n286) );
  INV_X1 U23 ( .A(n184), .ZN(n311) );
  INV_X1 U24 ( .A(n197), .ZN(n279) );
  INV_X1 U25 ( .A(n148), .ZN(n308) );
  INV_X1 U26 ( .A(n73), .ZN(n296) );
  INV_X1 U27 ( .A(n218), .ZN(n313) );
  INV_X1 U28 ( .A(n199), .ZN(n280) );
  INV_X1 U29 ( .A(n170), .ZN(n329) );
  INV_X1 U30 ( .A(n124), .ZN(n312) );
  INV_X1 U31 ( .A(n81), .ZN(n325) );
  INV_X1 U32 ( .A(n195), .ZN(n319) );
  INV_X1 U33 ( .A(n67), .ZN(n276) );
  INV_X1 U34 ( .A(n158), .ZN(n302) );
  INV_X1 U35 ( .A(n92), .ZN(n295) );
  INV_X1 U36 ( .A(n183), .ZN(n320) );
  INV_X1 U37 ( .A(n84), .ZN(n314) );
  INV_X1 U38 ( .A(n146), .ZN(n310) );
  INV_X1 U39 ( .A(n108), .ZN(n303) );
  INV_X1 U40 ( .A(n91), .ZN(n306) );
  INV_X1 U41 ( .A(n97), .ZN(n305) );
  INV_X1 U42 ( .A(n153), .ZN(n317) );
  INV_X1 U43 ( .A(n79), .ZN(n326) );
  INV_X1 U45 ( .A(n193), .ZN(n331) );
  INV_X1 U46 ( .A(n163), .ZN(n283) );
  INV_X1 U48 ( .A(n151), .ZN(n318) );
  INV_X1 U49 ( .A(n99), .ZN(n288) );
  INV_X1 U50 ( .A(n211), .ZN(n285) );
  INV_X1 U51 ( .A(n89), .ZN(n298) );
  INV_X1 U52 ( .A(n98), .ZN(n289) );
  INV_X1 U53 ( .A(n196), .ZN(n291) );
  INV_X1 U54 ( .A(n229), .ZN(n277) );
  INV_X1 U55 ( .A(IR_IN_27), .ZN(n307) );
  INV_X1 U56 ( .A(IR_IN_28), .ZN(n304) );
  INV_X1 U57 ( .A(n135), .ZN(n332) );
  INV_X1 U58 ( .A(IR_IN_31), .ZN(n282) );
  INV_X1 U59 ( .A(IR_IN[5]), .ZN(n322) );
  INV_X1 U60 ( .A(IR_IN_30), .ZN(n297) );
  INV_X1 U61 ( .A(cw[2]), .ZN(n284) );
  INV_X1 U62 ( .A(IR_IN_29), .ZN(n299) );
  INV_X1 U64 ( .A(IR_IN_26), .ZN(n309) );
  INV_X1 U65 ( .A(IR_IN[3]), .ZN(n324) );
  INV_X1 U66 ( .A(IR_IN[0]), .ZN(n333) );
  INV_X1 U268 ( .A(IR_IN[2]), .ZN(n328) );
  INV_X1 U269 ( .A(n200), .ZN(n281) );
  INV_X1 U270 ( .A(IR_IN[4]), .ZN(n323) );
  DFFR_X1 \cw3_reg[13]  ( .D(cw2[13]), .CK(Clk), .RN(Rst), .Q(MUXA_SEL) );
  DFFR_X1 \cw2_reg[13]  ( .D(cw1[13]), .CK(Clk), .RN(Rst), .Q(cw2[13]) );
  DFFR_X1 \cw3_reg[12]  ( .D(cw2[12]), .CK(Clk), .RN(Rst), .Q(MUXB_SEL) );
  DFFR_X1 \cw1_reg[19]  ( .D(1'b1), .CK(Clk), .RN(Rst), .Q(IF_LATCH_EN) );
  DFFR_X1 \cw1_reg[18]  ( .D(1'b1), .CK(Clk), .RN(Rst), .Q(cw1[18]) );
  SDFFR_X1 \cw1_reg[17]  ( .D(n286), .SI(1'b0), .SE(n327), .CK(Clk), .RN(Rst), 
        .Q(cw1[17]) );
  DFFR_X1 \cw1_reg[16]  ( .D(n252), .CK(Clk), .RN(Rst), .Q(cw1[16]) );
  DFFR_X1 \cw1_reg[15]  ( .D(cw[15]), .CK(Clk), .RN(Rst), .Q(cw1[15]) );
  DFFR_X1 \cw1_reg[14]  ( .D(cw[14]), .CK(Clk), .RN(Rst), .Q(cw1[14]) );
  DFFR_X1 \cw1_reg[13]  ( .D(cw[13]), .CK(Clk), .RN(Rst), .Q(cw1[13]) );
  DFFR_X1 \cw1_reg[12]  ( .D(cw[12]), .CK(Clk), .RN(Rst), .Q(cw1[12]) );
  DFFR_X1 \cw1_reg[11]  ( .D(1'b1), .CK(Clk), .RN(Rst), .Q(cw1[11]) );
  DFFR_X1 \cw1_reg[10]  ( .D(n291), .CK(Clk), .RN(Rst), .Q(cw1[10]) );
  DFFR_X1 \cw1_reg[9]  ( .D(cw[9]), .CK(Clk), .RN(Rst), .Q(cw1[9]) );
  DFFR_X1 \cw1_reg[8]  ( .D(1'b1), .CK(Clk), .RN(Rst), .Q(cw1[8]) );
  DFFR_X1 \cw1_reg[7]  ( .D(n280), .CK(Clk), .RN(Rst), .Q(cw1[7]) );
  DFFR_X1 \cw1_reg[6]  ( .D(cw[6]), .CK(Clk), .RN(Rst), .Q(cw1[6]) );
  DFFR_X1 \cw1_reg[5]  ( .D(n281), .CK(Clk), .RN(Rst), .Q(cw1[5]) );
  DFFR_X1 \cw1_reg[4]  ( .D(cw[4]), .CK(Clk), .RN(Rst), .Q(cw1[4]) );
  DFFR_X1 \cw1_reg[3]  ( .D(cw[3]), .CK(Clk), .RN(Rst), .Q(cw1[3]) );
  DFFR_X1 \cw1_reg[2]  ( .D(cw[2]), .CK(Clk), .RN(Rst), .Q(cw1[2]) );
  SDFFR_X1 \cw1_reg[1]  ( .D(IR_IN_28), .SI(1'b0), .SE(n254), .CK(Clk), .RN(
        Rst), .Q(cw1[1]) );
  DFFR_X1 \cw1_reg[0]  ( .D(n337), .CK(Clk), .RN(Rst), .Q(cw1[0]) );
  DFFR_X1 \cw2_reg[18]  ( .D(cw1[18]), .CK(Clk), .RN(Rst), .Q(DEC_OUTREG_EN)
         );
  DFFR_X1 \cw2_reg[17]  ( .D(cw1[17]), .CK(Clk), .RN(Rst), .Q(IS_I_TYPE) );
  DFFR_X1 \cw2_reg[16]  ( .D(cw1[16]), .CK(Clk), .RN(Rst), .Q(RD1_EN) );
  DFFR_X1 \cw2_reg[15]  ( .D(cw1[15]), .CK(Clk), .RN(Rst), .Q(RD2_EN) );
  DFFR_X1 \cw2_reg[14]  ( .D(cw1[14]), .CK(Clk), .RN(Rst), .Q(ZERO_PADDING2)
         );
  DFFR_X1 \cw2_reg[12]  ( .D(cw1[12]), .CK(Clk), .RN(Rst), .Q(cw2[12]) );
  DFFR_X1 \cw2_reg[11]  ( .D(cw1[11]), .CK(Clk), .RN(Rst), .Q(cw2[11]) );
  DFFR_X1 \cw2_reg[10]  ( .D(cw1[10]), .CK(Clk), .RN(Rst), .Q(cw2[10]) );
  DFFR_X1 \cw2_reg[9]  ( .D(cw1[9]), .CK(Clk), .RN(Rst), .Q(cw2[9]) );
  DFFR_X1 \cw2_reg[8]  ( .D(cw1[8]), .CK(Clk), .RN(Rst), .Q(cw2[8]) );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(Clk), .RN(Rst), .Q(cw2[7]) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(Clk), .RN(Rst), .Q(cw2[6]) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(Clk), .RN(Rst), .Q(cw2[5]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(Clk), .RN(Rst), .Q(cw2[4]) );
  DFFR_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(Clk), .RN(Rst), .Q(cw2[3]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(Clk), .RN(Rst), .Q(cw2[2]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(Clk), .RN(Rst), .Q(cw2[1]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(Clk), .RN(Rst), .Q(cw2[0]) );
  DFFR_X1 \cw3_reg[11]  ( .D(cw2[11]), .CK(Clk), .RN(Rst), .Q(EXE_OUTREG_EN)
         );
  DFFR_X1 \cw3_reg[10]  ( .D(cw2[10]), .CK(Clk), .RN(Rst), .Q(EQ_COND) );
  DFFR_X1 \cw3_reg[9]  ( .D(cw2[9]), .CK(Clk), .RN(Rst), .Q(JUMP_EN) );
  DFFR_X1 \cw3_reg[8]  ( .D(cw2[8]), .CK(Clk), .RN(Rst), .Q(cw3[8]) );
  DFFR_X1 \cw3_reg[7]  ( .D(cw2[7]), .CK(Clk), .RN(Rst), .Q(cw3[7]) );
  DFFR_X1 \cw3_reg[6]  ( .D(cw2[6]), .CK(Clk), .RN(Rst), .Q(cw3[6]) );
  DFFR_X1 \cw3_reg[5]  ( .D(cw2[5]), .CK(Clk), .RN(Rst), .Q(cw3[5]) );
  DFFR_X1 \cw3_reg[4]  ( .D(cw2[4]), .CK(Clk), .RN(Rst), .Q(cw3[4]) );
  DFFR_X1 \cw3_reg[3]  ( .D(cw2[3]), .CK(Clk), .RN(Rst), .Q(cw3[3]) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .CK(Clk), .RN(Rst), .Q(cw3[2]) );
  DFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .CK(Clk), .RN(Rst), .Q(cw3[1]) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .CK(Clk), .RN(Rst), .Q(cw3[0]) );
  DFFR_X1 \cw4_reg[8]  ( .D(cw3[8]), .CK(Clk), .RN(Rst), .Q(MEM_OUTREG_EN) );
  DFFR_X1 \cw4_reg[7]  ( .D(cw3[7]), .CK(Clk), .RN(Rst), .Q(DRAM_WE) );
  DFFR_X1 \cw4_reg[6]  ( .D(cw3[6]), .CK(Clk), .RN(Rst), .Q(BYTE_LEN[1]) );
  DFFR_X1 \cw4_reg[5]  ( .D(cw3[5]), .CK(Clk), .RN(Rst), .Q(BYTE_LEN[0]) );
  DFFR_X1 \cw4_reg[4]  ( .D(cw3[4]), .CK(Clk), .RN(Rst), .Q(cw4[4]) );
  DFFR_X1 \cw4_reg[3]  ( .D(cw3[3]), .CK(Clk), .RN(Rst), .Q(cw4[3]) );
  DFFR_X1 \cw4_reg[2]  ( .D(cw3[2]), .CK(Clk), .RN(Rst), .Q(cw4[2]) );
  DFFR_X1 \cw4_reg[1]  ( .D(cw3[1]), .CK(Clk), .RN(Rst), .Q(cw4[1]) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3[0]), .CK(Clk), .RN(Rst), .Q(cw4[0]) );
  DFFR_X1 \cw5_reg[5]  ( .D(cw4[4]), .CK(Clk), .RN(Rst), .Q(WB_MUX_SEL[1]) );
  DFFR_X1 \cw5_reg[4]  ( .D(cw4[3]), .CK(Clk), .RN(Rst), .Q(WB_MUX_SEL[0]) );
  DFFR_X1 \cw5_reg[3]  ( .D(cw4[2]), .CK(Clk), .RN(Rst), .Q(JAL_REG31) );
  DFFR_X1 \cw5_reg[2]  ( .D(BYTE_LEN[0]), .CK(Clk), .RN(Rst), .Q(WB_CTRL_SIGN)
         );
  DFFR_X1 \cw5_reg[1]  ( .D(cw4[1]), .CK(Clk), .RN(Rst), .Q(ZERO_PADDING5) );
  DFFR_X1 \cw5_reg[0]  ( .D(cw4[0]), .CK(Clk), .RN(Rst), .Q(WR_EN) );
  DFFS_X1 \ALU_op1_reg[6]  ( .D(n38), .CK(Clk), .SN(Rst), .Q(ALU_op1[6]) );
  DFFR_X1 \ALU_op1_reg[5]  ( .D(\ALU_op[5] ), .CK(Clk), .RN(Rst), .Q(
        ALU_op1[5]) );
  DFFR_X1 \ALU_op1_reg[4]  ( .D(n63), .CK(Clk), .RN(Rst), .Q(ALU_op1[4]) );
  DFFS_X1 \ALU_op1_reg[3]  ( .D(n57), .CK(Clk), .SN(Rst), .Q(ALU_op1[3]) );
  DFFR_X1 \ALU_op1_reg[2]  ( .D(n336), .CK(Clk), .RN(Rst), .Q(ALU_op1[2]) );
  DFFS_X1 \ALU_op1_reg[1]  ( .D(n82), .CK(Clk), .SN(Rst), .Q(ALU_op1[1]) );
  DFFS_X1 \ALU_op1_reg[0]  ( .D(n46), .CK(Clk), .SN(Rst), .Q(ALU_op1[0]) );
  DFFR_X1 \ALU_op2_reg[5]  ( .D(ALU_op1[5]), .CK(Clk), .RN(Rst), .Q(ALU_op2[5]) );
  DFFR_X1 \ALU_op2_reg[4]  ( .D(ALU_op1[4]), .CK(Clk), .RN(Rst), .Q(ALU_op2[4]) );
  DFFR_X1 \ALU_op2_reg[2]  ( .D(ALU_op1[2]), .CK(Clk), .RN(Rst), .Q(ALU_op2[2]) );
  DFFR_X1 \ALU_op3_reg[5]  ( .D(ALU_op2[5]), .CK(Clk), .RN(Rst), .Q(
        \ALU_OPCODE[5] ) );
  DFFR_X1 \ALU_op3_reg[4]  ( .D(ALU_op2[4]), .CK(Clk), .RN(Rst), .Q(
        \ALU_OPCODE[4] ) );
  DFFR_X1 \ALU_op3_reg[2]  ( .D(ALU_op2[2]), .CK(Clk), .RN(Rst), .Q(
        \ALU_OPCODE[2] ) );
  DFFS_X1 \FPU_op1_reg[4]  ( .D(n26), .CK(Clk), .SN(Rst), .Q(FPU_op1[4]) );
  SDFFS_X1 \FPU_op1_reg[3]  ( .D(1'b1), .SI(IR_IN[3]), .SE(n253), .CK(Clk), 
        .SN(Rst), .Q(FPU_op1[3]) );
  SDFFS_X1 \FPU_op1_reg[2]  ( .D(1'b1), .SI(IR_IN[2]), .SE(n253), .CK(Clk), 
        .SN(Rst), .Q(FPU_op1[2]) );
  SDFFS_X1 \FPU_op1_reg[1]  ( .D(1'b1), .SI(IR_IN[1]), .SE(n253), .CK(Clk), 
        .SN(Rst), .Q(FPU_op1[1]) );
  SDFFR_X1 \FPU_op1_reg[0]  ( .D(IR_IN[0]), .SI(1'b0), .SE(n315), .CK(Clk), 
        .RN(Rst), .Q(FPU_op1[0]) );
  DFFR_X1 \FPU_op2_reg[0]  ( .D(FPU_op1[0]), .CK(Clk), .RN(Rst), .Q(FPU_op2[0]) );
  DFFR_X1 \FPU_op3_reg[0]  ( .D(FPU_op2[0]), .CK(Clk), .RN(Rst), .Q(
        FPU_OPCODE[0]) );
  DFFS_X1 \FPU_op2_reg[3]  ( .D(FPU_op1[3]), .CK(Clk), .SN(Rst), .Q(FPU_op2[3]) );
  DFFS_X1 \FPU_op2_reg[2]  ( .D(FPU_op1[2]), .CK(Clk), .SN(Rst), .Q(FPU_op2[2]) );
  DFFS_X1 \FPU_op2_reg[1]  ( .D(FPU_op1[1]), .CK(Clk), .SN(Rst), .Q(FPU_op2[1]) );
  DFFS_X1 \FPU_op2_reg[4]  ( .D(FPU_op1[4]), .CK(Clk), .SN(Rst), .Q(FPU_op2[4]) );
  DFFS_X1 \ALU_op3_reg[1]  ( .D(ALU_op2[1]), .CK(Clk), .SN(Rst), .Q(
        ALU_OPCODE[1]) );
  DFFS_X1 \ALU_op2_reg[1]  ( .D(ALU_op1[1]), .CK(Clk), .SN(Rst), .Q(ALU_op2[1]) );
  DFFS_X1 \FPU_op3_reg[4]  ( .D(FPU_op2[4]), .CK(Clk), .SN(Rst), .Q(
        FPU_OPCODE[4]) );
  DFFS_X1 \FPU_op3_reg[3]  ( .D(FPU_op2[3]), .CK(Clk), .SN(Rst), .Q(
        FPU_OPCODE[3]) );
  DFFS_X1 \FPU_op3_reg[2]  ( .D(FPU_op2[2]), .CK(Clk), .SN(Rst), .Q(
        FPU_OPCODE[2]) );
  DFFS_X1 \FPU_op3_reg[1]  ( .D(FPU_op2[1]), .CK(Clk), .SN(Rst), .Q(
        FPU_OPCODE[1]) );
  DFFS_X1 \ALU_op2_reg[6]  ( .D(ALU_op1[6]), .CK(Clk), .SN(Rst), .Q(ALU_op2[6]) );
  DFFS_X1 \ALU_op2_reg[3]  ( .D(ALU_op1[3]), .CK(Clk), .SN(Rst), .Q(ALU_op2[3]) );
  DFFS_X1 \ALU_op2_reg[0]  ( .D(ALU_op1[0]), .CK(Clk), .SN(Rst), .Q(ALU_op2[0]) );
  DFFS_X1 \ALU_op3_reg[6]  ( .D(ALU_op2[6]), .CK(Clk), .SN(Rst), .Q(
        ALU_OPCODE[6]) );
  DFFS_X1 \ALU_op3_reg[3]  ( .D(ALU_op2[3]), .CK(Clk), .SN(Rst), .Q(
        ALU_OPCODE[3]) );
  DFFS_X1 \ALU_op3_reg[0]  ( .D(ALU_op2[0]), .CK(Clk), .SN(Rst), .Q(
        ALU_OPCODE[0]) );
  OR4_X1 U9 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .A3(IR_IN[7]), .A4(IR_IN[10]), 
        .ZN(n334) );
  OR3_X1 U10 ( .A1(n172), .A2(n153), .A3(n76), .ZN(n335) );
  OR4_X1 U11 ( .A1(n118), .A2(n119), .A3(n279), .A4(n120), .ZN(n336) );
  OR4_X1 U12 ( .A1(n203), .A2(n293), .A3(n227), .A4(n217), .ZN(n337) );
  AND2_X1 U44 ( .A1(n173), .A2(n170), .ZN(n180) );
  AND2_X1 U47 ( .A1(n308), .A2(n83), .ZN(n74) );
  AND2_X1 U63 ( .A1(n26), .A2(n192), .ZN(n315) );
  AND2_X1 U76 ( .A1(IR_IN_26), .A2(n66), .ZN(n227) );
endmodule


module DLX ( Clock, ResetN, Instr_In, ProgCount_Out, DataMem_WrEn, 
        DataMem_BLen, DataMem_Addr, DataMem_Write, DataMem_Read );
  input [31:0] Instr_In;
  output [31:0] ProgCount_Out;
  output [1:0] DataMem_BLen;
  output [31:0] DataMem_Addr;
  output [31:0] DataMem_Write;
  input [31:0] DataMem_Read;
  input Clock, ResetN;
  output DataMem_WrEn;
  wire   IF_LATCH_EN, DEC_OUTREG_EN, IS_I_TYPE, RD1_EN, RD2_EN, WR_EN,
         JAL_REG31, ZERO_PADDING2, MUXA_SEL, MUXB_SEL, EXE_OUTREG_EN, EQ_COND,
         JUMP_EN, MEM_OUTREG_EN, DRAM_WE_INT, WB_CTRL_SIGN, ZERO_PADDING5;
  wire   [6:0] ALU_OPCODE;
  wire   [1:0] BYTE_LEN_INT;
  wire   [1:0] WB_MUX_SEL;
  wire   [31:0] IR_IN;

  DP_N_BITS_DATA32_N_BYTES_INST4_RF_ADDR5_N_BITS_JUMP26_N_BITS_IMM16 DATAPATH ( 
        .CLK(Clock), .RST(ResetN), .IF_LATCH_EN(IF_LATCH_EN), .DEC_OUTREG_EN(
        DEC_OUTREG_EN), .IS_I_TYPE(IS_I_TYPE), .RD1_EN(RD1_EN), .RD2_EN(RD2_EN), .WR_EN(WR_EN), .JAL_REG31(JAL_REG31), .ZERO_PADDING2(ZERO_PADDING2), 
        .MUXA_SEL(MUXA_SEL), .MUXB_SEL(MUXB_SEL), .EXE_OUTREG_EN(EXE_OUTREG_EN), .EQ_COND(EQ_COND), .JUMP_EN(JUMP_EN), .ALU_OPCODE(ALU_OPCODE), 
        .MEM_OUTREG_EN(MEM_OUTREG_EN), .BYTE_LEN_IN(BYTE_LEN_INT), .DRAM_WE(
        DRAM_WE_INT), .DRAM_WE_OUT(DataMem_WrEn), .BYTE_LEN_OUT(DataMem_BLen), 
        .WB_MUX_SEL(WB_MUX_SEL), .WB_CTRL_SIGN(WB_CTRL_SIGN), .ZERO_PADDING5(
        ZERO_PADDING5), .IR_IN(IR_IN), .PC_OUT(ProgCount_Out), 
        .MEM_DATA_OUT_INT(DataMem_Read), .MEM_ADDR_OUT(DataMem_Addr), 
        .MEM_DATA_IN_PRIME(DataMem_Write) );
  CU_HW_MICRO_SIZE154_FUNC_SIZE11_OPCODE_SIZE6_IR_SIZE32_CW_SIZE20 CONTROL ( 
        .Clk(Clock), .Rst(ResetN), .IR_IN(Instr_In), .IF_LATCH_EN(IF_LATCH_EN), 
        .DEC_OUTREG_EN(DEC_OUTREG_EN), .IS_I_TYPE(IS_I_TYPE), .RD1_EN(RD1_EN), 
        .RD2_EN(RD2_EN), .ZERO_PADDING2(ZERO_PADDING2), .MUXA_SEL(MUXA_SEL), 
        .MUXB_SEL(MUXB_SEL), .EXE_OUTREG_EN(EXE_OUTREG_EN), .EQ_COND(EQ_COND), 
        .JUMP_EN(JUMP_EN), .ALU_OPCODE(ALU_OPCODE), .MEM_OUTREG_EN(
        MEM_OUTREG_EN), .DRAM_WE(DRAM_WE_INT), .BYTE_LEN(BYTE_LEN_INT), 
        .WB_MUX_SEL(WB_MUX_SEL), .JAL_REG31(JAL_REG31), .WB_CTRL_SIGN(
        WB_CTRL_SIGN), .ZERO_PADDING5(ZERO_PADDING5), .WR_EN(WR_EN) );
  DFFR_X1 \IR_IN_reg[31]  ( .D(Instr_In[31]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[31]) );
  DFFR_X1 \IR_IN_reg[30]  ( .D(Instr_In[30]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[30]) );
  DFFR_X1 \IR_IN_reg[29]  ( .D(Instr_In[29]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[29]) );
  DFFR_X1 \IR_IN_reg[28]  ( .D(Instr_In[28]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[28]) );
  DFFR_X1 \IR_IN_reg[27]  ( .D(Instr_In[27]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[27]) );
  DFFR_X1 \IR_IN_reg[26]  ( .D(Instr_In[26]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[26]) );
  DFFR_X1 \IR_IN_reg[25]  ( .D(Instr_In[25]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[25]) );
  DFFR_X1 \IR_IN_reg[24]  ( .D(Instr_In[24]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[24]) );
  DFFR_X1 \IR_IN_reg[23]  ( .D(Instr_In[23]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[23]) );
  DFFR_X1 \IR_IN_reg[22]  ( .D(Instr_In[22]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[22]) );
  DFFR_X1 \IR_IN_reg[21]  ( .D(Instr_In[21]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[21]) );
  DFFR_X1 \IR_IN_reg[20]  ( .D(Instr_In[20]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[20]) );
  DFFR_X1 \IR_IN_reg[19]  ( .D(Instr_In[19]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[19]) );
  DFFR_X1 \IR_IN_reg[18]  ( .D(Instr_In[18]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[18]) );
  DFFR_X1 \IR_IN_reg[17]  ( .D(Instr_In[17]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[17]) );
  DFFR_X1 \IR_IN_reg[16]  ( .D(Instr_In[16]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[16]) );
  DFFR_X1 \IR_IN_reg[15]  ( .D(Instr_In[15]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[15]) );
  DFFR_X1 \IR_IN_reg[14]  ( .D(Instr_In[14]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[14]) );
  DFFR_X1 \IR_IN_reg[13]  ( .D(Instr_In[13]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[13]) );
  DFFR_X1 \IR_IN_reg[12]  ( .D(Instr_In[12]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[12]) );
  DFFR_X1 \IR_IN_reg[11]  ( .D(Instr_In[11]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[11]) );
  DFFR_X1 \IR_IN_reg[10]  ( .D(Instr_In[10]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[10]) );
  DFFR_X1 \IR_IN_reg[9]  ( .D(Instr_In[9]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[9]) );
  DFFR_X1 \IR_IN_reg[8]  ( .D(Instr_In[8]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[8]) );
  DFFR_X1 \IR_IN_reg[7]  ( .D(Instr_In[7]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[7]) );
  DFFR_X1 \IR_IN_reg[6]  ( .D(Instr_In[6]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[6]) );
  DFFR_X1 \IR_IN_reg[5]  ( .D(Instr_In[5]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[5]) );
  DFFR_X1 \IR_IN_reg[4]  ( .D(Instr_In[4]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[4]) );
  DFFR_X1 \IR_IN_reg[3]  ( .D(Instr_In[3]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[3]) );
  DFFR_X1 \IR_IN_reg[2]  ( .D(Instr_In[2]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[2]) );
  DFFR_X1 \IR_IN_reg[1]  ( .D(Instr_In[1]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[1]) );
  DFFR_X1 \IR_IN_reg[0]  ( .D(Instr_In[0]), .CK(Clock), .RN(ResetN), .Q(
        IR_IN[0]) );
endmodule

